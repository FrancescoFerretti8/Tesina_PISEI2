magic
tech sky130A
magscale 1 2
timestamp 1750758279
<< viali >>
rect -636 -6664 -564 -6492
rect -342 -6662 -270 -6490
rect -66 -6660 6 -6488
rect 228 -6662 300 -6490
rect 482 -6664 554 -6492
rect 772 -6666 844 -6494
<< metal1 >>
rect 5254 1225 5454 1230
rect -1202 1007 1916 1207
rect 4754 1025 5454 1225
rect 5254 976 5454 1025
rect 5254 770 5454 776
rect -1200 597 -1000 598
rect -1200 595 1666 597
rect -1200 398 1892 595
rect 4764 421 6404 621
rect -1098 397 1892 398
rect 1542 395 1892 397
rect -1198 -285 1894 -85
rect 4812 -230 5958 -30
rect 5758 -548 5958 -230
rect 5752 -748 5758 -548
rect 5958 -748 5964 -548
rect 5248 -1282 5254 -1082
rect 5454 -1282 5460 -1082
rect 5254 -1583 5454 -1282
rect -1218 -1801 1934 -1601
rect 4772 -1783 5454 -1583
rect 1708 -1802 1774 -1801
rect 5254 -1838 5454 -1783
rect 5254 -2044 5454 -2038
rect 6204 -2187 6404 421
rect -1212 -2406 1770 -2206
rect 4770 -2387 6404 -2187
rect 1542 -2408 1762 -2406
rect 5758 -2578 5958 -2572
rect 5758 -2837 5958 -2778
rect 1668 -2893 1836 -2892
rect -1192 -3093 1912 -2893
rect 4788 -3037 5958 -2837
rect 5758 -3232 5958 -3037
rect -262 -3524 -256 -3324
rect -56 -3524 -50 -3324
rect 5752 -3432 5758 -3232
rect 5958 -3432 5964 -3232
rect -256 -3774 -56 -3524
rect 6204 -3688 6404 -2387
rect -532 -4224 220 -3774
rect 596 -3898 1276 -3842
rect 6204 -3888 6846 -3688
rect 596 -4098 4910 -3898
rect 596 -4154 1276 -4098
rect 1218 -4399 1798 -4392
rect 4710 -4399 4910 -4098
rect 5248 -4236 5254 -4036
rect 5454 -4236 5460 -4036
rect 5254 -4399 5454 -4236
rect -1260 -4612 1798 -4399
rect 4652 -4599 5454 -4399
rect -1260 -4614 1285 -4612
rect 5254 -4620 5454 -4599
rect 5254 -4826 5454 -4820
rect 6204 -5003 6404 -3888
rect 1260 -5229 1266 -5029
rect 1466 -5229 1836 -5029
rect 4708 -5203 6404 -5003
rect 5758 -5442 5958 -5436
rect 5758 -5653 5958 -5642
rect -1258 -5710 1435 -5703
rect -1258 -5910 1792 -5710
rect 4706 -5853 5958 -5653
rect -1258 -5918 1435 -5910
rect -730 -6488 4886 -6476
rect 5758 -6478 5958 -5853
rect -730 -6490 -66 -6488
rect -730 -6492 -342 -6490
rect -730 -6664 -636 -6492
rect -564 -6662 -342 -6492
rect -270 -6660 -66 -6490
rect 6 -6490 4886 -6488
rect 6 -6660 228 -6490
rect -270 -6662 228 -6660
rect 300 -6492 4886 -6490
rect 300 -6662 482 -6492
rect -564 -6664 482 -6662
rect 554 -6494 4886 -6492
rect 554 -6664 772 -6494
rect -730 -6666 772 -6664
rect 844 -6666 4886 -6494
rect -730 -6676 4886 -6666
rect 4686 -7081 4886 -6676
rect 5752 -6678 5758 -6478
rect 5958 -6678 5964 -6478
rect 5248 -6878 5254 -6678
rect 5454 -6878 5460 -6678
rect 5254 -7081 5454 -6878
rect -1246 -7308 1788 -7108
rect 4660 -7281 5458 -7081
rect 6204 -7685 6404 -5203
rect 808 -7911 1812 -7711
rect 4684 -7800 6404 -7685
rect 4684 -7885 6402 -7800
rect -1242 -8586 -1018 -8386
rect -818 -8586 -812 -8386
rect -559 -9118 -333 -8319
rect 58 -8544 734 -8372
rect 808 -8544 1008 -7911
rect 5758 -7976 5958 -7970
rect 5758 -8335 5958 -8176
rect 58 -8744 1008 -8544
rect 1116 -8386 1316 -8380
rect 1316 -8586 1728 -8386
rect 4690 -8535 5958 -8335
rect 1116 -8592 1316 -8586
rect 58 -8860 734 -8744
rect 5758 -9118 5958 -8535
rect -559 -9318 5958 -9118
rect -559 -9331 -333 -9318
<< via1 >>
rect 5254 776 5454 976
rect 5758 -748 5958 -548
rect 5254 -1282 5454 -1082
rect 5254 -2038 5454 -1838
rect 5758 -2778 5958 -2578
rect -256 -3524 -56 -3324
rect 5758 -3432 5958 -3232
rect 5254 -4236 5454 -4036
rect 5254 -4820 5454 -4620
rect 1266 -5229 1466 -5029
rect 5758 -5642 5958 -5442
rect 5758 -6678 5958 -6478
rect 5254 -6878 5454 -6678
rect -1018 -8586 -818 -8386
rect 5758 -8176 5958 -7976
rect 1116 -8586 1316 -8386
<< metal2 >>
rect 5248 776 5254 976
rect 5454 776 5460 976
rect 5254 -1082 5454 776
rect 5254 -1288 5454 -1282
rect 5758 -548 5958 -542
rect 5248 -2038 5254 -1838
rect 5454 -2038 5460 -1838
rect -256 -3324 -56 -3318
rect -56 -3524 1466 -3324
rect -256 -3530 -56 -3524
rect 1266 -5029 1466 -3524
rect 5254 -4036 5454 -2038
rect 5758 -2578 5958 -748
rect 5752 -2778 5758 -2578
rect 5958 -2778 5964 -2578
rect 5254 -4242 5454 -4236
rect 5758 -3232 5958 -3226
rect 5248 -4820 5254 -4620
rect 5454 -4820 5460 -4620
rect 1266 -5235 1466 -5229
rect 5254 -6678 5454 -4820
rect 5758 -5442 5958 -3432
rect 5752 -5642 5758 -5442
rect 5958 -5642 5964 -5442
rect 5254 -6884 5454 -6878
rect 5758 -6478 5958 -6472
rect 5758 -7976 5958 -6678
rect 5752 -8176 5758 -7976
rect 5958 -8176 5964 -7976
rect -1018 -8386 -818 -8380
rect -818 -8586 1116 -8386
rect 1316 -8586 1322 -8386
rect -1018 -8592 -818 -8586
use pass_gate  x1
timestamp 1750758113
transform 1 0 1274 0 1 165
box 418 -835 3696 1565
use pass_gate  x2
timestamp 1750758113
transform 1 0 1292 0 1 -2643
box 418 -835 3696 1565
use pass_gate  x3
timestamp 1750758113
transform 1 0 1218 0 1 -5459
box 418 -835 3696 1565
use pass_gate  x4
timestamp 1750758113
transform 1 0 1194 0 1 -8141
box 418 -835 3696 1565
use sky130_fd_pr__res_high_po_0p35_B5WUZC  XR1
timestamp 1750754129
transform 1 0 117 0 1 -6324
box -201 -2682 201 2682
use sky130_fd_pr__res_high_po_0p35_B5WUZC  XR2
timestamp 1750754129
transform 1 0 663 0 1 -6350
box -201 -2682 201 2682
use sky130_fd_pr__res_high_po_0p35_B5WUZC  XR3
timestamp 1750754129
transform 1 0 -459 0 1 -6318
box -201 -2682 201 2682
<< labels >>
flabel metal1 6646 -3888 6846 -3688 0 FreeSans 256 0 0 0 out
port 8 nsew
flabel metal1 -1212 -2406 -1012 -2206 0 FreeSans 256 0 0 0 A1
port 6 nsew
flabel metal1 -1200 398 -1000 598 0 FreeSans 256 0 0 0 A0
port 3 nsew
flabel metal1 -1202 1007 1916 1207 0 FreeSans 256 0 0 0 n0
port 24 nsew
flabel metal1 -1198 -285 -998 -85 0 FreeSans 256 0 0 0 p0
port 26 nsew
flabel metal1 -1218 -1801 -1018 -1601 0 FreeSans 256 0 0 0 n1
port 28 nsew
flabel metal1 -1192 -3093 -992 -2893 0 FreeSans 256 0 0 0 p1
port 30 nsew
flabel metal1 -1248 -4602 -1042 -4402 0 FreeSans 256 0 0 0 n2
port 34 nsew
flabel metal1 -1250 -5910 -1030 -5710 0 FreeSans 256 0 0 0 p2
port 35 nsew
flabel metal1 -1246 -7308 -910 -7108 0 FreeSans 256 0 0 0 n3
port 37 nsew
flabel metal1 -1242 -8586 -1018 -8386 0 FreeSans 256 0 0 0 p3
port 39 nsew
flabel metal1 5254 976 5454 1230 0 FreeSans 256 0 0 0 VSS
port 41 nsew
flabel metal1 5758 -9318 5958 -8176 0 FreeSans 256 0 0 0 VDD
port 43 nsew
<< end >>
