** sch_path: /home/ttuser/Progetto_PISEI/xschem/pass_gate.sch
.subckt pass_gate VDD VSS pin Ain uscita nin
*.PININFO Ain:I pin:I nin:I VDD:I VSS:I uscita:O
XM2 Ain nin uscita VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=8 nf=8 m=1
XM3 uscita pin Ain VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=16 nf=16 m=1
.ends
.end
