magic
tech sky130A
magscale 1 2
timestamp 1750763685
<< metal1 >>
rect 7232 44498 7238 44558
rect 7298 44498 7304 44558
rect 17406 44552 17412 44612
rect 17472 44552 17478 44612
rect 6852 44052 7052 44058
rect 7238 44052 7298 44498
rect 8888 44372 8894 44432
rect 8954 44372 8960 44432
rect 7784 44176 7790 44236
rect 7850 44176 7856 44236
rect 7790 44052 7850 44176
rect 8336 44150 8342 44210
rect 8402 44150 8408 44210
rect 8342 44052 8402 44150
rect 8894 44052 8954 44372
rect 10544 44360 10550 44420
rect 10610 44360 10616 44420
rect 11648 44372 11654 44432
rect 11714 44372 11720 44432
rect 9446 44352 9506 44358
rect 9446 44052 9506 44292
rect 9992 44134 9998 44194
rect 10058 44134 10064 44194
rect 9998 44052 10058 44134
rect 10550 44052 10610 44360
rect 11096 44240 11102 44300
rect 11162 44240 11168 44300
rect 11102 44052 11162 44240
rect 11654 44052 11714 44372
rect 16970 44052 17170 44058
rect 17412 44052 17472 44552
rect 18824 44388 18830 44448
rect 18890 44388 18896 44448
rect 19376 44436 19382 44496
rect 19442 44436 19448 44496
rect 17720 44282 17726 44342
rect 17786 44282 17792 44342
rect 17726 44052 17786 44282
rect 18272 44102 18278 44162
rect 18338 44102 18344 44162
rect 18278 44052 18338 44102
rect 18830 44052 18890 44388
rect 19382 44052 19442 44436
rect 20480 44342 20486 44402
rect 20546 44342 20552 44402
rect 22136 44348 22142 44408
rect 22202 44348 22208 44408
rect 27668 44360 27724 44366
rect 19928 44232 19934 44292
rect 19994 44232 20000 44292
rect 19934 44052 19994 44232
rect 20486 44052 20546 44342
rect 21032 44288 21038 44348
rect 21098 44288 21104 44348
rect 21038 44052 21098 44288
rect 21584 44276 21590 44336
rect 21650 44276 21656 44336
rect 21590 44052 21650 44276
rect 22142 44052 22202 44348
rect 22688 44278 22694 44338
rect 22754 44278 22760 44338
rect 23240 44286 23246 44346
rect 23306 44286 23312 44346
rect 22694 44052 22754 44278
rect 23246 44052 23306 44286
rect 27126 44162 27182 44168
rect 7052 43852 12048 44052
rect 12248 43852 12254 44052
rect 17170 43852 23390 44052
rect 23590 43852 23596 44052
rect 6852 43846 7052 43852
rect 16970 43846 17170 43852
rect 27126 42776 27182 44106
rect 27120 42720 27126 42776
rect 27182 42720 27188 42776
rect 11512 41710 11568 41716
rect 22394 41710 22450 41716
rect 27668 41710 27724 44304
rect 11568 41654 16670 41710
rect 16726 41654 16732 41710
rect 22450 41654 27724 41710
rect 11512 41648 11568 41654
rect 22394 41648 22450 41654
rect 6180 39872 6236 39878
rect 6180 35206 6236 39816
rect 21226 39472 21282 39478
rect 27126 39472 27182 39478
rect 11148 39416 11864 39472
rect 11920 39416 11926 39472
rect 21282 39416 27126 39472
rect 6174 35150 6180 35206
rect 6236 35150 6242 35206
rect 11148 35020 11204 39416
rect 21226 39410 21282 39416
rect 27126 39410 27182 39416
rect 11142 34964 11148 35020
rect 11204 34964 11210 35020
rect 27572 28430 27772 28436
rect 27572 28224 27772 28230
rect 20120 27660 20240 27666
rect 20240 27540 20634 27660
rect 20120 27534 20240 27540
rect 12932 26328 12988 26334
rect 12988 26272 20780 26328
rect 12932 26266 12988 26272
rect 20032 24996 20152 25002
rect 20152 24876 20798 24996
rect 20032 24870 20152 24876
rect 13854 23562 21066 23618
rect 13854 16138 13910 23562
rect 28462 22800 30522 23000
rect 19760 22192 19880 22198
rect 19880 22072 20870 22192
rect 19760 22066 19880 22072
rect 20182 21318 20188 21518
rect 20388 21318 20872 21518
rect 14706 20786 20780 20842
rect 13848 16082 13854 16138
rect 13910 16082 13916 16138
rect 14706 16028 14762 20786
rect 19870 19326 19990 19332
rect 19990 19206 20704 19326
rect 19870 19200 19990 19206
rect 19454 18714 19654 18720
rect 19654 18514 20826 18714
rect 19454 18508 19654 18514
rect 16188 18008 21000 18064
rect 14700 15972 14706 16028
rect 14762 15972 14768 16028
rect 16188 16008 16244 18008
rect 18776 17754 18782 17954
rect 18982 17754 18988 17954
rect 16182 15952 16188 16008
rect 16244 15952 16250 16008
rect 18782 13016 18982 17754
rect 27080 17258 27280 18090
rect 27080 17052 27280 17058
rect 22544 13016 22744 13022
rect 18782 12816 22544 13016
rect 22544 12810 22744 12816
rect 30322 1688 30522 22800
rect 30322 1660 30542 1688
rect 30362 1052 30542 1660
rect 30356 872 30362 1052
rect 30542 872 30548 1052
<< via1 >>
rect 7238 44498 7298 44558
rect 17412 44552 17472 44612
rect 8894 44372 8954 44432
rect 7790 44176 7850 44236
rect 8342 44150 8402 44210
rect 10550 44360 10610 44420
rect 11654 44372 11714 44432
rect 9446 44292 9506 44352
rect 9998 44134 10058 44194
rect 11102 44240 11162 44300
rect 18830 44388 18890 44448
rect 19382 44436 19442 44496
rect 17726 44282 17786 44342
rect 18278 44102 18338 44162
rect 20486 44342 20546 44402
rect 22142 44348 22202 44408
rect 19934 44232 19994 44292
rect 21038 44288 21098 44348
rect 21590 44276 21650 44336
rect 22694 44278 22754 44338
rect 23246 44286 23306 44346
rect 27668 44304 27724 44360
rect 27126 44106 27182 44162
rect 6852 43852 7052 44052
rect 12048 43852 12248 44052
rect 16970 43852 17170 44052
rect 23390 43852 23590 44052
rect 27126 42720 27182 42776
rect 11512 41654 11568 41710
rect 16670 41654 16726 41710
rect 22394 41654 22450 41710
rect 6180 39816 6236 39872
rect 11864 39416 11920 39472
rect 21226 39416 21282 39472
rect 27126 39416 27182 39472
rect 6180 35150 6236 35206
rect 11148 34964 11204 35020
rect 27572 28230 27772 28430
rect 20120 27540 20240 27660
rect 12932 26272 12988 26328
rect 20032 24876 20152 24996
rect 19760 22072 19880 22192
rect 20188 21318 20388 21518
rect 13854 16082 13910 16138
rect 19870 19206 19990 19326
rect 19454 18514 19654 18714
rect 14706 15972 14762 16028
rect 18782 17754 18982 17954
rect 16188 15952 16244 16008
rect 27080 17058 27280 17258
rect 22544 12816 22744 13016
rect 30362 872 30542 1052
<< metal2 >>
rect 22694 44784 22754 44786
rect 7238 44762 7298 44764
rect 12758 44762 12818 44764
rect 6686 44710 6746 44712
rect 6679 44654 6688 44710
rect 6744 44654 6753 44710
rect 7231 44706 7240 44762
rect 7296 44706 7305 44762
rect 12751 44706 12760 44762
rect 12816 44706 12825 44762
rect 22142 44734 22202 44736
rect 6134 44376 6194 44378
rect 6127 44320 6136 44376
rect 6192 44320 6201 44376
rect 3763 44052 3953 44056
rect 6134 44052 6194 44320
rect 6686 44052 6746 44654
rect 7238 44558 7298 44706
rect 10550 44684 10610 44686
rect 8894 44668 8954 44670
rect 7790 44630 7850 44632
rect 7783 44574 7792 44630
rect 7848 44574 7857 44630
rect 8887 44612 8896 44668
rect 8952 44612 8961 44668
rect 10543 44628 10552 44684
rect 10608 44628 10617 44684
rect 11102 44662 11162 44664
rect 7238 44492 7298 44498
rect 7790 44236 7850 44574
rect 8342 44550 8402 44552
rect 8335 44494 8344 44550
rect 8400 44494 8409 44550
rect 7790 44170 7850 44176
rect 8342 44210 8402 44494
rect 8894 44432 8954 44612
rect 9446 44598 9506 44600
rect 9998 44598 10058 44600
rect 9439 44542 9448 44598
rect 9504 44542 9513 44598
rect 9991 44542 10000 44598
rect 10056 44542 10065 44598
rect 8894 44366 8954 44372
rect 9446 44352 9506 44542
rect 9440 44292 9446 44352
rect 9506 44292 9512 44352
rect 8342 44144 8402 44150
rect 9998 44194 10058 44542
rect 10550 44420 10610 44628
rect 11095 44606 11104 44662
rect 11160 44606 11169 44662
rect 11656 44616 11712 44623
rect 11654 44614 11714 44616
rect 10550 44354 10610 44360
rect 11102 44300 11162 44606
rect 11654 44558 11656 44614
rect 11712 44558 11714 44614
rect 11654 44432 11714 44558
rect 12206 44550 12266 44552
rect 12199 44494 12208 44550
rect 12264 44494 12273 44550
rect 11654 44366 11714 44372
rect 12206 44342 12266 44494
rect 12206 44282 12482 44342
rect 11102 44234 11162 44240
rect 9998 44128 10058 44134
rect 12048 44052 12248 44058
rect 12422 44052 12482 44282
rect 12758 44052 12818 44706
rect 20486 44686 20546 44688
rect 18830 44684 18890 44686
rect 13310 44630 13370 44632
rect 17726 44630 17786 44632
rect 13303 44574 13312 44630
rect 13368 44574 13377 44630
rect 17176 44612 17232 44619
rect 17412 44612 17472 44618
rect 17174 44610 17412 44612
rect 14414 44604 14474 44606
rect 13310 44052 13370 44574
rect 14407 44548 14416 44604
rect 14472 44548 14481 44604
rect 17174 44554 17176 44610
rect 17232 44554 17412 44610
rect 17174 44552 17412 44554
rect 17719 44574 17728 44630
rect 17784 44574 17793 44630
rect 18823 44628 18832 44684
rect 18888 44628 18897 44684
rect 19382 44666 19442 44668
rect 18278 44604 18338 44606
rect 16622 44550 16682 44552
rect 13862 44466 13922 44468
rect 13855 44410 13864 44466
rect 13920 44410 13929 44466
rect 13862 44052 13922 44410
rect 14414 44052 14474 44548
rect 14966 44536 15026 44538
rect 14959 44480 14968 44536
rect 15024 44480 15033 44536
rect 15518 44498 15578 44500
rect 14966 44052 15026 44480
rect 15511 44442 15520 44498
rect 15576 44442 15585 44498
rect 16615 44494 16624 44550
rect 16680 44494 16689 44550
rect 17176 44545 17232 44552
rect 17412 44546 17472 44552
rect 15518 44052 15578 44442
rect 16070 44360 16130 44362
rect 16063 44304 16072 44360
rect 16128 44304 16137 44360
rect 16070 44052 16130 44304
rect 16622 44052 16682 44494
rect 17726 44342 17786 44574
rect 18271 44548 18280 44604
rect 18336 44548 18345 44604
rect 17726 44276 17786 44282
rect 18278 44162 18338 44548
rect 18830 44448 18890 44628
rect 19375 44610 19384 44666
rect 19440 44610 19449 44666
rect 19934 44642 19994 44644
rect 19382 44496 19442 44610
rect 19927 44586 19936 44642
rect 19992 44586 20001 44642
rect 20479 44630 20488 44686
rect 20544 44630 20553 44686
rect 21590 44678 21650 44680
rect 22135 44678 22144 44734
rect 22200 44678 22209 44734
rect 22687 44728 22696 44784
rect 22752 44728 22761 44784
rect 19382 44430 19442 44436
rect 18830 44382 18890 44388
rect 19934 44292 19994 44586
rect 20486 44402 20546 44630
rect 21583 44622 21592 44678
rect 21648 44622 21657 44678
rect 21038 44592 21098 44594
rect 21031 44536 21040 44592
rect 21096 44536 21105 44592
rect 20486 44336 20546 44342
rect 21038 44348 21098 44536
rect 21038 44282 21098 44288
rect 21590 44336 21650 44622
rect 22142 44408 22202 44678
rect 22142 44342 22202 44348
rect 21590 44270 21650 44276
rect 22694 44338 22754 44728
rect 28214 44664 28274 44666
rect 23246 44650 23306 44652
rect 23239 44594 23248 44650
rect 23304 44594 23313 44650
rect 28207 44608 28216 44664
rect 28272 44608 28281 44664
rect 28766 44654 28826 44656
rect 23246 44346 23306 44594
rect 27666 44584 27726 44593
rect 27666 44515 27726 44524
rect 27124 44504 27184 44513
rect 27124 44435 27184 44444
rect 23246 44280 23306 44286
rect 22694 44272 22754 44278
rect 19934 44226 19994 44232
rect 27126 44162 27182 44435
rect 27668 44360 27724 44515
rect 27662 44304 27668 44360
rect 27724 44304 27730 44360
rect 27120 44106 27126 44162
rect 27182 44106 27188 44162
rect 18278 44096 18338 44102
rect 23390 44052 23590 44058
rect 28214 44052 28274 44608
rect 28759 44598 28768 44654
rect 28824 44598 28833 44654
rect 28766 44052 28826 44598
rect 3758 44047 6852 44052
rect 3758 43857 3763 44047
rect 3953 43857 6852 44047
rect 3758 43852 6852 43857
rect 7052 43852 7058 44052
rect 12248 43852 16970 44052
rect 17170 43852 17176 44052
rect 23590 43852 29394 44052
rect 3763 43848 3953 43852
rect 12048 43846 12248 43852
rect 23390 43846 23590 43852
rect 27126 42776 27182 42782
rect 16670 41710 16726 41716
rect 6180 41654 11512 41710
rect 11568 41654 11574 41710
rect 16726 41654 22394 41710
rect 22450 41654 22456 41710
rect 6180 39872 6236 41654
rect 16670 41648 16726 41654
rect 6174 39816 6180 39872
rect 6236 39816 6242 39872
rect 11864 39472 11920 39478
rect 27126 39472 27182 42720
rect 11920 39416 21226 39472
rect 21282 39416 21288 39472
rect 27120 39416 27126 39472
rect 27182 39416 27188 39472
rect 11864 39410 11920 39416
rect 6180 35206 6236 35212
rect 6180 31264 6236 35150
rect 11148 35020 11204 35026
rect 11148 31264 11204 34964
rect 15017 29908 15026 30308
rect 15426 29908 28794 30308
rect 13563 29048 13673 29052
rect 13558 29043 19934 29048
rect 13558 28933 13563 29043
rect 13673 28933 19934 29043
rect 13558 28928 19934 28933
rect 13563 28924 13673 28928
rect 19814 27660 19934 28928
rect 27572 28430 27772 29908
rect 27566 28230 27572 28430
rect 27772 28230 27778 28430
rect 19814 27540 20120 27660
rect 20240 27540 20246 27660
rect 12926 26272 12932 26328
rect 12988 26272 12994 26328
rect 4892 12170 4948 15376
rect 7376 13206 7432 15398
rect 9860 14198 9916 15394
rect 12344 15204 12400 15376
rect 12932 15204 12988 26272
rect 13563 25240 13673 25244
rect 13558 25235 20152 25240
rect 13558 25125 13563 25235
rect 13673 25125 20152 25235
rect 13558 25120 20152 25125
rect 13563 25116 13673 25120
rect 20032 24996 20152 25120
rect 20026 24876 20032 24996
rect 20152 24876 20158 24996
rect 19754 22072 19760 22192
rect 19880 22072 19886 22192
rect 13563 21432 13673 21436
rect 19760 21432 19880 22072
rect 13558 21427 19880 21432
rect 13558 21317 13563 21427
rect 13673 21317 19880 21427
rect 13558 21312 19880 21317
rect 20188 21518 20388 21524
rect 13563 21308 13673 21312
rect 19864 19206 19870 19326
rect 19990 19206 19996 19326
rect 18782 18514 19454 18714
rect 19654 18514 19660 18714
rect 18782 17954 18982 18514
rect 18782 17748 18982 17754
rect 13561 17624 13671 17628
rect 19870 17624 19990 19206
rect 13556 17619 19990 17624
rect 13556 17509 13561 17619
rect 13671 17509 19990 17619
rect 13556 17504 19990 17509
rect 13561 17500 13671 17504
rect 12344 15148 12988 15204
rect 13854 16138 13910 16144
rect 13854 14198 13910 16082
rect 20188 16088 20388 21318
rect 27074 17058 27080 17258
rect 27280 17058 27286 17258
rect 9860 14142 13910 14198
rect 14706 16028 14762 16034
rect 14706 13206 14762 15972
rect 7376 13150 14762 13206
rect 16188 16008 16244 16014
rect 16188 12170 16244 15952
rect 20188 15888 25728 16088
rect 22538 12816 22544 13016
rect 22744 12816 22750 13016
rect 4892 12114 16244 12170
rect 22544 7802 22744 12816
rect 22544 7593 22744 7602
rect 25528 3556 25728 15888
rect 27080 14600 27280 17058
rect 27080 14391 27280 14400
rect 26474 3556 26674 3565
rect 25528 3356 26474 3556
rect 26474 3347 26674 3356
rect 30362 1052 30542 1058
rect 30362 593 30542 872
rect 30358 423 30367 593
rect 30537 423 30546 593
rect 30362 418 30542 423
<< via2 >>
rect 6688 44654 6744 44710
rect 7240 44706 7296 44762
rect 12760 44706 12816 44762
rect 6136 44320 6192 44376
rect 7792 44574 7848 44630
rect 8896 44612 8952 44668
rect 10552 44628 10608 44684
rect 8344 44494 8400 44550
rect 9448 44542 9504 44598
rect 10000 44542 10056 44598
rect 11104 44606 11160 44662
rect 11656 44558 11712 44614
rect 12208 44494 12264 44550
rect 13312 44574 13368 44630
rect 14416 44548 14472 44604
rect 17176 44554 17232 44610
rect 17728 44574 17784 44630
rect 18832 44628 18888 44684
rect 13864 44410 13920 44466
rect 14968 44480 15024 44536
rect 15520 44442 15576 44498
rect 16624 44494 16680 44550
rect 16072 44304 16128 44360
rect 18280 44548 18336 44604
rect 19384 44610 19440 44666
rect 19936 44586 19992 44642
rect 20488 44630 20544 44686
rect 22144 44678 22200 44734
rect 22696 44728 22752 44784
rect 21592 44622 21648 44678
rect 21040 44536 21096 44592
rect 23248 44594 23304 44650
rect 28216 44608 28272 44664
rect 27666 44524 27726 44584
rect 27124 44444 27184 44504
rect 28768 44598 28824 44654
rect 3763 43857 3953 44047
rect 15026 29908 15426 30308
rect 13563 28933 13673 29043
rect 13563 25125 13673 25235
rect 13563 21317 13673 21427
rect 13561 17509 13671 17619
rect 22544 7602 22744 7802
rect 27080 14400 27280 14600
rect 26474 3356 26674 3556
rect 30367 423 30537 593
<< metal3 >>
rect 6678 44950 6684 45014
rect 6748 44950 6754 45014
rect 7230 44962 7236 45026
rect 7300 44962 7306 45026
rect 7782 44962 7788 45026
rect 7852 44962 7858 45026
rect 6686 44715 6746 44950
rect 7238 44767 7298 44962
rect 7235 44762 7301 44767
rect 6683 44710 6749 44715
rect 6126 44618 6132 44682
rect 6196 44618 6202 44682
rect 6683 44654 6688 44710
rect 6744 44654 6749 44710
rect 7235 44706 7240 44762
rect 7296 44706 7301 44762
rect 7235 44701 7301 44706
rect 6683 44649 6749 44654
rect 7790 44635 7850 44962
rect 8334 44950 8340 45014
rect 8404 44950 8410 45014
rect 8886 44968 8892 45032
rect 8956 44968 8962 45032
rect 7787 44630 7853 44635
rect 6134 44381 6194 44618
rect 7787 44574 7792 44630
rect 7848 44574 7853 44630
rect 7787 44569 7853 44574
rect 8342 44555 8402 44950
rect 8894 44673 8954 44968
rect 9438 44952 9444 45016
rect 9508 44952 9514 45016
rect 9990 44968 9996 45032
rect 10060 44968 10066 45032
rect 8891 44668 8957 44673
rect 8891 44612 8896 44668
rect 8952 44612 8957 44668
rect 8891 44607 8957 44612
rect 9446 44603 9506 44952
rect 9998 44603 10058 44968
rect 10542 44950 10548 45014
rect 10612 44950 10618 45014
rect 11094 44950 11100 45014
rect 11164 44950 11170 45014
rect 11646 44950 11652 45014
rect 11716 44950 11722 45014
rect 12198 44978 12204 45042
rect 12268 44978 12274 45042
rect 10550 44689 10610 44950
rect 10547 44684 10613 44689
rect 10547 44628 10552 44684
rect 10608 44628 10613 44684
rect 11102 44667 11162 44950
rect 10547 44623 10613 44628
rect 11099 44662 11165 44667
rect 11099 44606 11104 44662
rect 11160 44606 11165 44662
rect 11654 44619 11714 44950
rect 9443 44598 9509 44603
rect 8339 44550 8405 44555
rect 8339 44494 8344 44550
rect 8400 44494 8405 44550
rect 9443 44542 9448 44598
rect 9504 44542 9509 44598
rect 9443 44537 9509 44542
rect 9995 44598 10061 44603
rect 11099 44601 11165 44606
rect 11651 44614 11717 44619
rect 9995 44542 10000 44598
rect 10056 44542 10061 44598
rect 11651 44558 11656 44614
rect 11712 44558 11717 44614
rect 11651 44553 11717 44558
rect 12206 44555 12266 44978
rect 12750 44950 12756 45014
rect 12820 44950 12826 45014
rect 13302 44968 13308 45032
rect 13372 44968 13378 45032
rect 12758 44767 12818 44950
rect 12755 44762 12821 44767
rect 12755 44706 12760 44762
rect 12816 44706 12821 44762
rect 12755 44701 12821 44706
rect 13310 44635 13370 44968
rect 13854 44962 13860 45026
rect 13924 44962 13930 45026
rect 14406 44968 14412 45032
rect 14476 44968 14482 45032
rect 14958 44968 14964 45032
rect 15028 44968 15034 45032
rect 16068 45014 16132 45020
rect 13307 44630 13373 44635
rect 13307 44574 13312 44630
rect 13368 44574 13373 44630
rect 13307 44569 13373 44574
rect 9995 44537 10061 44542
rect 12203 44550 12269 44555
rect 8339 44489 8405 44494
rect 12203 44494 12208 44550
rect 12264 44494 12269 44550
rect 12203 44489 12269 44494
rect 13862 44471 13922 44962
rect 14414 44609 14474 44968
rect 14411 44604 14477 44609
rect 14411 44548 14416 44604
rect 14472 44548 14477 44604
rect 14411 44543 14477 44548
rect 14966 44541 15026 44968
rect 15510 44950 15516 45014
rect 15580 44950 15586 45014
rect 16062 44950 16068 45014
rect 16132 44950 16138 45014
rect 16614 44950 16620 45014
rect 16684 44950 16690 45014
rect 17166 44950 17172 45014
rect 17236 44950 17242 45014
rect 17718 44978 17724 45042
rect 17788 44978 17794 45042
rect 14963 44536 15029 44541
rect 14963 44480 14968 44536
rect 15024 44480 15029 44536
rect 15518 44503 15578 44950
rect 16068 44944 16132 44950
rect 14963 44475 15029 44480
rect 15515 44498 15581 44503
rect 13859 44466 13925 44471
rect 13859 44410 13864 44466
rect 13920 44410 13925 44466
rect 15515 44442 15520 44498
rect 15576 44442 15581 44498
rect 15515 44437 15581 44442
rect 13859 44405 13925 44410
rect 6131 44376 6197 44381
rect 6131 44320 6136 44376
rect 6192 44320 6197 44376
rect 16070 44365 16130 44944
rect 16622 44555 16682 44950
rect 17174 44615 17234 44950
rect 17726 44635 17786 44978
rect 18270 44952 18276 45016
rect 18340 44952 18346 45016
rect 18822 44952 18828 45016
rect 18892 44952 18898 45016
rect 17723 44630 17789 44635
rect 17171 44610 17237 44615
rect 16619 44550 16685 44555
rect 16619 44494 16624 44550
rect 16680 44494 16685 44550
rect 17171 44554 17176 44610
rect 17232 44554 17237 44610
rect 17723 44574 17728 44630
rect 17784 44574 17789 44630
rect 18278 44609 18338 44952
rect 18830 44689 18890 44952
rect 19374 44950 19380 45014
rect 19444 44950 19450 45014
rect 19926 44950 19932 45014
rect 19996 44950 20002 45014
rect 20478 44950 20484 45014
rect 20548 44950 20554 45014
rect 21030 44954 21036 45018
rect 21100 44954 21106 45018
rect 18827 44684 18893 44689
rect 18827 44628 18832 44684
rect 18888 44628 18893 44684
rect 19382 44671 19442 44950
rect 18827 44623 18893 44628
rect 19379 44666 19445 44671
rect 19379 44610 19384 44666
rect 19440 44610 19445 44666
rect 19934 44647 19994 44950
rect 20486 44691 20546 44950
rect 20483 44686 20549 44691
rect 17723 44569 17789 44574
rect 18275 44604 18341 44609
rect 19379 44605 19445 44610
rect 19931 44642 19997 44647
rect 17171 44549 17237 44554
rect 18275 44548 18280 44604
rect 18336 44548 18341 44604
rect 19931 44586 19936 44642
rect 19992 44586 19997 44642
rect 20483 44630 20488 44686
rect 20544 44630 20549 44686
rect 20483 44625 20549 44630
rect 21038 44597 21098 44954
rect 21582 44950 21588 45014
rect 21652 44950 21658 45014
rect 22134 44950 22140 45014
rect 22204 44950 22210 45014
rect 22686 44986 22692 45050
rect 22756 44986 22762 45050
rect 21590 44683 21650 44950
rect 22142 44739 22202 44950
rect 22694 44789 22754 44986
rect 23238 44950 23244 45014
rect 23308 44950 23314 45014
rect 28206 44956 28212 45020
rect 28276 44956 28282 45020
rect 22691 44784 22757 44789
rect 22139 44734 22205 44739
rect 21587 44678 21653 44683
rect 21587 44622 21592 44678
rect 21648 44622 21653 44678
rect 22139 44678 22144 44734
rect 22200 44678 22205 44734
rect 22691 44728 22696 44784
rect 22752 44728 22757 44784
rect 22691 44723 22757 44728
rect 22139 44673 22205 44678
rect 23246 44655 23306 44950
rect 27664 44750 27728 44756
rect 21587 44617 21653 44622
rect 23243 44650 23309 44655
rect 19931 44581 19997 44586
rect 21035 44592 21101 44597
rect 18275 44543 18341 44548
rect 21035 44536 21040 44592
rect 21096 44536 21101 44592
rect 23243 44594 23248 44650
rect 23304 44594 23309 44650
rect 27096 44628 27102 44692
rect 27166 44690 27172 44692
rect 27166 44630 27198 44690
rect 27664 44680 27728 44686
rect 27166 44628 27184 44630
rect 23243 44589 23309 44594
rect 21035 44531 21101 44536
rect 27124 44509 27184 44628
rect 27666 44589 27726 44680
rect 28214 44669 28274 44956
rect 28758 44950 28764 45014
rect 28828 44950 28834 45014
rect 28211 44664 28277 44669
rect 28211 44608 28216 44664
rect 28272 44608 28277 44664
rect 28766 44659 28826 44950
rect 28211 44603 28277 44608
rect 28763 44654 28829 44659
rect 28763 44598 28768 44654
rect 28824 44598 28829 44654
rect 28763 44593 28829 44598
rect 27661 44584 27731 44589
rect 27661 44524 27666 44584
rect 27726 44524 27731 44584
rect 27661 44519 27731 44524
rect 16619 44489 16685 44494
rect 27119 44504 27189 44509
rect 27119 44444 27124 44504
rect 27184 44444 27189 44504
rect 27119 44439 27189 44444
rect 6131 44315 6197 44320
rect 16067 44360 16133 44365
rect 16067 44304 16072 44360
rect 16128 44304 16133 44360
rect 16067 44299 16133 44304
rect 1001 44151 1199 44157
rect 1000 43852 1001 44052
rect 1199 44047 3958 44052
rect 1199 43857 3763 44047
rect 3953 43857 3958 44047
rect 1199 43852 3958 43857
rect 1001 43747 1199 43753
rect 2265 30308 2663 30313
rect 15021 30308 15431 30313
rect 210 29908 216 30308
rect 616 30307 2664 30308
rect 616 29909 2265 30307
rect 2663 29909 2664 30307
rect 616 29908 2664 29909
rect 13440 29908 13446 30308
rect 13846 29908 15026 30308
rect 15426 29908 15431 30308
rect 2265 29903 2663 29908
rect 15021 29903 15431 29908
rect 13558 29043 13678 29048
rect 13558 28933 13563 29043
rect 13673 28933 13678 29043
rect 13558 28928 13678 28933
rect 13558 25235 13678 25240
rect 13558 25125 13563 25235
rect 13673 25125 13678 25235
rect 13558 25120 13678 25125
rect 13558 21427 13678 21432
rect 13558 21317 13563 21427
rect 13673 21317 13678 21427
rect 13558 21312 13678 21317
rect 13556 17619 13676 17624
rect 13556 17509 13561 17619
rect 13671 17509 13676 17619
rect 13556 17504 13676 17509
rect 27075 14600 27285 14605
rect 27075 14400 27080 14600
rect 27280 14400 27285 14600
rect 27075 14395 27285 14400
rect 17403 13692 17677 13697
rect 27080 13692 27280 14395
rect 17402 13691 27394 13692
rect 17402 13417 17403 13691
rect 17677 13417 27394 13691
rect 17402 13416 27394 13417
rect 17403 13411 17677 13416
rect 22539 7802 22749 7807
rect 22539 7602 22544 7802
rect 22744 7602 22749 7802
rect 22539 7597 22749 7602
rect 22544 5428 22744 7597
rect 22544 5222 22744 5228
rect 26469 3556 26679 3561
rect 26469 3356 26474 3556
rect 26674 3356 26679 3556
rect 26469 3351 26679 3356
rect 26474 1518 26674 3351
rect 26474 1312 26674 1318
rect 30362 593 30542 598
rect 30362 423 30367 593
rect 30537 423 30542 593
rect 30362 199 30542 423
rect 30357 21 30363 199
rect 30541 21 30547 199
rect 30362 20 30542 21
<< via3 >>
rect 6684 44950 6748 45014
rect 7236 44962 7300 45026
rect 7788 44962 7852 45026
rect 6132 44618 6196 44682
rect 8340 44950 8404 45014
rect 8892 44968 8956 45032
rect 9444 44952 9508 45016
rect 9996 44968 10060 45032
rect 10548 44950 10612 45014
rect 11100 44950 11164 45014
rect 11652 44950 11716 45014
rect 12204 44978 12268 45042
rect 12756 44950 12820 45014
rect 13308 44968 13372 45032
rect 13860 44962 13924 45026
rect 14412 44968 14476 45032
rect 14964 44968 15028 45032
rect 15516 44950 15580 45014
rect 16068 44950 16132 45014
rect 16620 44950 16684 45014
rect 17172 44950 17236 45014
rect 17724 44978 17788 45042
rect 18276 44952 18340 45016
rect 18828 44952 18892 45016
rect 19380 44950 19444 45014
rect 19932 44950 19996 45014
rect 20484 44950 20548 45014
rect 21036 44954 21100 45018
rect 21588 44950 21652 45014
rect 22140 44950 22204 45014
rect 22692 44986 22756 45050
rect 23244 44950 23308 45014
rect 28212 44956 28276 45020
rect 27102 44628 27166 44692
rect 27664 44686 27728 44750
rect 28764 44950 28828 45014
rect 1001 43753 1199 44151
rect 216 29908 616 30308
rect 2265 29909 2663 30307
rect 13446 29908 13846 30308
rect 17403 13417 17677 13691
rect 22544 5228 22744 5428
rect 26474 1318 26674 1518
rect 30363 21 30541 199
<< metal4 >>
rect 6134 44683 6194 45152
rect 6686 45015 6746 45152
rect 7238 45027 7298 45152
rect 7790 45027 7850 45152
rect 7235 45026 7301 45027
rect 6683 45014 6749 45015
rect 6683 44950 6684 45014
rect 6748 44950 6749 45014
rect 7235 44962 7236 45026
rect 7300 44962 7301 45026
rect 7235 44961 7301 44962
rect 7787 45026 7853 45027
rect 7787 44962 7788 45026
rect 7852 44962 7853 45026
rect 8342 45015 8402 45152
rect 8894 45033 8954 45152
rect 8891 45032 8957 45033
rect 7787 44961 7853 44962
rect 8339 45014 8405 45015
rect 7238 44952 7298 44961
rect 7790 44952 7850 44961
rect 6683 44949 6749 44950
rect 8339 44950 8340 45014
rect 8404 44950 8405 45014
rect 8891 44968 8892 45032
rect 8956 44968 8957 45032
rect 9446 45017 9506 45152
rect 9998 45033 10058 45152
rect 9995 45032 10061 45033
rect 8891 44967 8957 44968
rect 9443 45016 9509 45017
rect 8894 44952 8954 44967
rect 9443 44952 9444 45016
rect 9508 44952 9509 45016
rect 9995 44968 9996 45032
rect 10060 44968 10061 45032
rect 10550 45015 10610 45152
rect 11102 45015 11162 45152
rect 11654 45015 11714 45152
rect 12206 45043 12266 45152
rect 12203 45042 12269 45043
rect 9995 44967 10061 44968
rect 10547 45014 10613 45015
rect 9998 44952 10058 44967
rect 9443 44951 9509 44952
rect 8339 44949 8405 44950
rect 10547 44950 10548 45014
rect 10612 44950 10613 45014
rect 10547 44949 10613 44950
rect 11099 45014 11165 45015
rect 11099 44950 11100 45014
rect 11164 44950 11165 45014
rect 11099 44949 11165 44950
rect 11651 45014 11717 45015
rect 11651 44950 11652 45014
rect 11716 44950 11717 45014
rect 12203 44978 12204 45042
rect 12268 44978 12269 45042
rect 12758 45015 12818 45152
rect 13310 45033 13370 45152
rect 13307 45032 13373 45033
rect 12203 44977 12269 44978
rect 12755 45014 12821 45015
rect 12206 44952 12266 44977
rect 11651 44949 11717 44950
rect 12755 44950 12756 45014
rect 12820 44950 12821 45014
rect 13307 44968 13308 45032
rect 13372 44968 13373 45032
rect 13862 45027 13922 45152
rect 14414 45033 14474 45152
rect 14966 45033 15026 45152
rect 14411 45032 14477 45033
rect 13307 44967 13373 44968
rect 13859 45026 13925 45027
rect 13310 44952 13370 44967
rect 13859 44962 13860 45026
rect 13924 44962 13925 45026
rect 14411 44968 14412 45032
rect 14476 44968 14477 45032
rect 14411 44967 14477 44968
rect 14963 45032 15029 45033
rect 14963 44968 14964 45032
rect 15028 44968 15029 45032
rect 15518 45015 15578 45152
rect 16070 45015 16130 45152
rect 16622 45015 16682 45152
rect 17174 45015 17234 45152
rect 17726 45043 17786 45152
rect 17723 45042 17789 45043
rect 14963 44967 15029 44968
rect 15515 45014 15581 45015
rect 13859 44961 13925 44962
rect 13862 44952 13922 44961
rect 14414 44952 14474 44967
rect 14966 44952 15026 44967
rect 12755 44949 12821 44950
rect 15515 44950 15516 45014
rect 15580 44950 15581 45014
rect 15515 44949 15581 44950
rect 16067 45014 16133 45015
rect 16067 44950 16068 45014
rect 16132 44950 16133 45014
rect 16067 44949 16133 44950
rect 16619 45014 16685 45015
rect 16619 44950 16620 45014
rect 16684 44950 16685 45014
rect 16619 44949 16685 44950
rect 17171 45014 17237 45015
rect 17171 44950 17172 45014
rect 17236 44950 17237 45014
rect 17723 44978 17724 45042
rect 17788 44978 17789 45042
rect 18278 45017 18338 45152
rect 18830 45017 18890 45152
rect 17723 44977 17789 44978
rect 18275 45016 18341 45017
rect 17726 44952 17786 44977
rect 18275 44952 18276 45016
rect 18340 44952 18341 45016
rect 18275 44951 18341 44952
rect 18827 45016 18893 45017
rect 18827 44952 18828 45016
rect 18892 44952 18893 45016
rect 19382 45015 19442 45152
rect 19934 45015 19994 45152
rect 20486 45015 20546 45152
rect 21038 45019 21098 45152
rect 21035 45018 21101 45019
rect 18827 44951 18893 44952
rect 19379 45014 19445 45015
rect 17171 44949 17237 44950
rect 19379 44950 19380 45014
rect 19444 44950 19445 45014
rect 19379 44949 19445 44950
rect 19931 45014 19997 45015
rect 19931 44950 19932 45014
rect 19996 44950 19997 45014
rect 19931 44949 19997 44950
rect 20483 45014 20549 45015
rect 20483 44950 20484 45014
rect 20548 44950 20549 45014
rect 21035 44954 21036 45018
rect 21100 44954 21101 45018
rect 21590 45015 21650 45152
rect 22142 45015 22202 45152
rect 22694 45051 22754 45152
rect 22691 45050 22757 45051
rect 21035 44953 21101 44954
rect 21587 45014 21653 45015
rect 21038 44952 21098 44953
rect 20483 44949 20549 44950
rect 21587 44950 21588 45014
rect 21652 44950 21653 45014
rect 21587 44949 21653 44950
rect 22139 45014 22205 45015
rect 22139 44950 22140 45014
rect 22204 44950 22205 45014
rect 22691 44986 22692 45050
rect 22756 44986 22757 45050
rect 23246 45015 23306 45152
rect 22691 44985 22757 44986
rect 23243 45014 23309 45015
rect 22694 44952 22754 44985
rect 22139 44949 22205 44950
rect 23243 44950 23244 45014
rect 23308 44950 23309 45014
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 45006 27170 45152
rect 27104 44952 27170 45006
rect 27662 45008 27722 45152
rect 28214 45021 28274 45152
rect 28211 45020 28277 45021
rect 27662 44952 27726 45008
rect 28211 44956 28212 45020
rect 28276 44956 28277 45020
rect 28766 45015 28826 45152
rect 28211 44955 28277 44956
rect 28763 45014 28829 45015
rect 28214 44952 28274 44955
rect 23243 44949 23309 44950
rect 27104 44693 27164 44952
rect 27666 44751 27726 44952
rect 28763 44950 28764 45014
rect 28828 44950 28829 45014
rect 29318 44952 29378 45152
rect 28763 44949 28829 44950
rect 27663 44750 27729 44751
rect 27101 44692 27167 44693
rect 6131 44682 6197 44683
rect 6131 44618 6132 44682
rect 6196 44618 6197 44682
rect 27101 44628 27102 44692
rect 27166 44628 27167 44692
rect 27663 44686 27664 44750
rect 27728 44686 27729 44750
rect 27663 44685 27729 44686
rect 27101 44627 27167 44628
rect 6131 44617 6197 44618
rect 200 30309 600 44152
rect 800 44151 1200 44152
rect 800 43753 1001 44151
rect 1199 43753 1200 44151
rect 200 30308 617 30309
rect 200 29908 216 30308
rect 616 29908 617 30308
rect 200 29907 617 29908
rect 200 1000 600 29907
rect 800 13692 1200 43753
rect 13445 30308 13847 30309
rect 2264 30307 13446 30308
rect 2264 29909 2265 30307
rect 2663 29909 13446 30307
rect 2264 29908 13446 29909
rect 13846 29908 13847 30308
rect 6244 28888 6644 29908
rect 7710 28844 8110 29908
rect 9178 28788 9578 29908
rect 10632 28820 11032 29908
rect 13445 29907 13847 29908
rect 7032 13692 7308 17590
rect 8496 13692 8772 17542
rect 9984 13692 10260 17602
rect 11424 13692 11700 17660
rect 800 13691 17678 13692
rect 800 13417 17403 13691
rect 17677 13417 17678 13691
rect 800 13416 17678 13417
rect 800 1000 1200 13416
rect 22543 5428 22745 5429
rect 22543 5228 22544 5428
rect 22744 5228 22745 5428
rect 22543 5227 22745 5228
rect 22544 200 22744 5227
rect 26473 1518 26675 1519
rect 26473 1318 26474 1518
rect 26674 1318 26675 1518
rect 26473 1317 26675 1318
rect 26474 200 26674 1317
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22544 56 22814 200
rect 26474 162 26678 200
rect 22634 0 22814 56
rect 26498 0 26678 162
rect 30362 199 30542 200
rect 30362 21 30363 199
rect 30541 21 30542 199
rect 30362 0 30542 21
use Decoder  Decoder_0
timestamp 1750763685
transform 1 0 3678 0 1 15320
box 1210 0 10000 16000
use Mux  Mux_0
timestamp 1750758279
transform 1 0 21826 0 -1 19112
box -1260 -9331 6846 1730
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 800 28236 1200 28636 0 FreeSans 1600 0 0 0 VGND
port 54 nsew
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
