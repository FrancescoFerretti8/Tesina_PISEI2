magic
tech sky130A
magscale 1 2
timestamp 1750763685
<< error_p >>
rect 6837 13413 6871 13447
rect 2697 13277 2731 13311
rect 7481 13277 7515 13311
rect 2881 13209 2915 13243
rect 7021 13209 7055 13243
rect 7389 13141 7423 13175
rect 7297 12937 7331 12971
rect 7297 12801 7331 12835
rect 7481 12801 7515 12835
rect 7481 10625 7515 10659
rect 7297 10421 7331 10455
rect 7021 10217 7055 10251
rect 7389 10217 7423 10251
rect 6929 10013 6963 10047
rect 7297 9537 7331 9571
rect 7481 9401 7515 9435
rect 7113 6409 7147 6443
rect 6929 6273 6963 6307
rect 7297 6273 7331 6307
rect 7481 6069 7515 6103
rect 6929 5865 6963 5899
rect 7297 5865 7331 5899
rect 7389 5661 7423 5695
rect 3157 3077 3191 3111
rect 2789 3009 2823 3043
rect 2973 3009 3007 3043
rect 2973 2805 3007 2839
rect 2697 2397 2731 2431
rect 2329 2329 2363 2363
<< viali >>
rect 6837 13413 6871 13447
rect 2697 13277 2731 13311
rect 7481 13277 7515 13311
rect 2881 13209 2915 13243
rect 7021 13209 7055 13243
rect 7389 13141 7423 13175
rect 7297 12937 7331 12971
rect 7297 12801 7331 12835
rect 7481 12801 7515 12835
rect 7481 10625 7515 10659
rect 7297 10421 7331 10455
rect 7021 10217 7055 10251
rect 7389 10217 7423 10251
rect 6929 10013 6963 10047
rect 7297 9537 7331 9571
rect 7481 9401 7515 9435
rect 7113 6409 7147 6443
rect 6929 6273 6963 6307
rect 7297 6273 7331 6307
rect 7481 6069 7515 6103
rect 6929 5865 6963 5899
rect 7297 5865 7331 5899
rect 7389 5661 7423 5695
rect 7389 3485 7423 3519
rect 7205 3417 7239 3451
rect 7021 3349 7055 3383
rect 3157 3077 3191 3111
rect 2789 3009 2823 3043
rect 2973 3009 3007 3043
rect 3709 3009 3743 3043
rect 6101 3009 6135 3043
rect 6469 3009 6503 3043
rect 6929 3009 6963 3043
rect 7113 3009 7147 3043
rect 7481 3009 7515 3043
rect 3617 2941 3651 2975
rect 5549 2941 5583 2975
rect 6009 2941 6043 2975
rect 6745 2941 6779 2975
rect 3525 2873 3559 2907
rect 5917 2873 5951 2907
rect 6653 2873 6687 2907
rect 2973 2805 3007 2839
rect 3893 2805 3927 2839
rect 6285 2805 6319 2839
rect 7297 2805 7331 2839
rect 2697 2397 2731 2431
rect 3893 2397 3927 2431
rect 6193 2397 6227 2431
rect 7021 2397 7055 2431
rect 7297 2397 7331 2431
rect 2329 2329 2363 2363
rect 3985 2261 4019 2295
rect 6285 2261 6319 2295
rect 6929 2261 6963 2295
rect 7481 2261 7515 2295
<< metal1 >>
rect 2024 13626 7912 13648
rect 2024 13574 2606 13626
rect 2658 13574 2670 13626
rect 2722 13574 2734 13626
rect 2786 13574 2798 13626
rect 2850 13574 2862 13626
rect 2914 13574 4078 13626
rect 4130 13574 4142 13626
rect 4194 13574 4206 13626
rect 4258 13574 4270 13626
rect 4322 13574 4334 13626
rect 4386 13574 5550 13626
rect 5602 13574 5614 13626
rect 5666 13574 5678 13626
rect 5730 13574 5742 13626
rect 5794 13574 5806 13626
rect 5858 13574 7022 13626
rect 7074 13574 7086 13626
rect 7138 13574 7150 13626
rect 7202 13574 7214 13626
rect 7266 13574 7278 13626
rect 7330 13574 7912 13626
rect 2024 13552 7912 13574
rect 6825 13447 6883 13453
rect 6825 13413 6837 13447
rect 6871 13444 6883 13447
rect 8294 13444 8300 13456
rect 6871 13416 8300 13444
rect 6871 13413 6883 13416
rect 6825 13407 6883 13413
rect 8294 13404 8300 13416
rect 8352 13404 8358 13456
rect 2498 13268 2504 13320
rect 2556 13308 2562 13320
rect 2685 13311 2743 13317
rect 2685 13308 2697 13311
rect 2556 13280 2697 13308
rect 2556 13268 2562 13280
rect 2685 13277 2697 13280
rect 2731 13277 2743 13311
rect 2685 13271 2743 13277
rect 7466 13268 7472 13320
rect 7524 13268 7530 13320
rect 2869 13243 2927 13249
rect 2869 13209 2881 13243
rect 2915 13240 2927 13243
rect 6914 13240 6920 13252
rect 2915 13212 6920 13240
rect 2915 13209 2927 13212
rect 2869 13203 2927 13209
rect 6914 13200 6920 13212
rect 6972 13200 6978 13252
rect 7009 13243 7067 13249
rect 7009 13209 7021 13243
rect 7055 13240 7067 13243
rect 7282 13240 7288 13252
rect 7055 13212 7288 13240
rect 7055 13209 7067 13212
rect 7009 13203 7067 13209
rect 7282 13200 7288 13212
rect 7340 13200 7346 13252
rect 7377 13175 7435 13181
rect 7377 13141 7389 13175
rect 7423 13172 7435 13175
rect 7466 13172 7472 13184
rect 7423 13144 7472 13172
rect 7423 13141 7435 13144
rect 7377 13135 7435 13141
rect 7466 13132 7472 13144
rect 7524 13132 7530 13184
rect 2024 13082 8072 13104
rect 2024 13030 3342 13082
rect 3394 13030 3406 13082
rect 3458 13030 3470 13082
rect 3522 13030 3534 13082
rect 3586 13030 3598 13082
rect 3650 13030 4814 13082
rect 4866 13030 4878 13082
rect 4930 13030 4942 13082
rect 4994 13030 5006 13082
rect 5058 13030 5070 13082
rect 5122 13030 6286 13082
rect 6338 13030 6350 13082
rect 6402 13030 6414 13082
rect 6466 13030 6478 13082
rect 6530 13030 6542 13082
rect 6594 13030 7758 13082
rect 7810 13030 7822 13082
rect 7874 13030 7886 13082
rect 7938 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8072 13082
rect 2024 13008 8072 13030
rect 7282 12928 7288 12980
rect 7340 12928 7346 12980
rect 6914 12792 6920 12844
rect 6972 12832 6978 12844
rect 7285 12835 7343 12841
rect 7285 12832 7297 12835
rect 6972 12804 7297 12832
rect 6972 12792 6978 12804
rect 7285 12801 7297 12804
rect 7331 12801 7343 12835
rect 7285 12795 7343 12801
rect 7466 12792 7472 12844
rect 7524 12792 7530 12844
rect 2024 12538 7912 12560
rect 2024 12486 2606 12538
rect 2658 12486 2670 12538
rect 2722 12486 2734 12538
rect 2786 12486 2798 12538
rect 2850 12486 2862 12538
rect 2914 12486 4078 12538
rect 4130 12486 4142 12538
rect 4194 12486 4206 12538
rect 4258 12486 4270 12538
rect 4322 12486 4334 12538
rect 4386 12486 5550 12538
rect 5602 12486 5614 12538
rect 5666 12486 5678 12538
rect 5730 12486 5742 12538
rect 5794 12486 5806 12538
rect 5858 12486 7022 12538
rect 7074 12486 7086 12538
rect 7138 12486 7150 12538
rect 7202 12486 7214 12538
rect 7266 12486 7278 12538
rect 7330 12486 7912 12538
rect 2024 12464 7912 12486
rect 2024 11994 8072 12016
rect 2024 11942 3342 11994
rect 3394 11942 3406 11994
rect 3458 11942 3470 11994
rect 3522 11942 3534 11994
rect 3586 11942 3598 11994
rect 3650 11942 4814 11994
rect 4866 11942 4878 11994
rect 4930 11942 4942 11994
rect 4994 11942 5006 11994
rect 5058 11942 5070 11994
rect 5122 11942 6286 11994
rect 6338 11942 6350 11994
rect 6402 11942 6414 11994
rect 6466 11942 6478 11994
rect 6530 11942 6542 11994
rect 6594 11942 7758 11994
rect 7810 11942 7822 11994
rect 7874 11942 7886 11994
rect 7938 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8072 11994
rect 2024 11920 8072 11942
rect 2024 11450 7912 11472
rect 2024 11398 2606 11450
rect 2658 11398 2670 11450
rect 2722 11398 2734 11450
rect 2786 11398 2798 11450
rect 2850 11398 2862 11450
rect 2914 11398 4078 11450
rect 4130 11398 4142 11450
rect 4194 11398 4206 11450
rect 4258 11398 4270 11450
rect 4322 11398 4334 11450
rect 4386 11398 5550 11450
rect 5602 11398 5614 11450
rect 5666 11398 5678 11450
rect 5730 11398 5742 11450
rect 5794 11398 5806 11450
rect 5858 11398 7022 11450
rect 7074 11398 7086 11450
rect 7138 11398 7150 11450
rect 7202 11398 7214 11450
rect 7266 11398 7278 11450
rect 7330 11398 7912 11450
rect 2024 11376 7912 11398
rect 2024 10906 8072 10928
rect 2024 10854 3342 10906
rect 3394 10854 3406 10906
rect 3458 10854 3470 10906
rect 3522 10854 3534 10906
rect 3586 10854 3598 10906
rect 3650 10854 4814 10906
rect 4866 10854 4878 10906
rect 4930 10854 4942 10906
rect 4994 10854 5006 10906
rect 5058 10854 5070 10906
rect 5122 10854 6286 10906
rect 6338 10854 6350 10906
rect 6402 10854 6414 10906
rect 6466 10854 6478 10906
rect 6530 10854 6542 10906
rect 6594 10854 7758 10906
rect 7810 10854 7822 10906
rect 7874 10854 7886 10906
rect 7938 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8072 10906
rect 2024 10832 8072 10854
rect 7374 10616 7380 10668
rect 7432 10656 7438 10668
rect 7469 10659 7527 10665
rect 7469 10656 7481 10659
rect 7432 10628 7481 10656
rect 7432 10616 7438 10628
rect 7469 10625 7481 10628
rect 7515 10625 7527 10659
rect 7469 10619 7527 10625
rect 7285 10455 7343 10461
rect 7285 10421 7297 10455
rect 7331 10452 7343 10455
rect 7558 10452 7564 10464
rect 7331 10424 7564 10452
rect 7331 10421 7343 10424
rect 7285 10415 7343 10421
rect 7558 10412 7564 10424
rect 7616 10412 7622 10464
rect 2024 10362 7912 10384
rect 2024 10310 2606 10362
rect 2658 10310 2670 10362
rect 2722 10310 2734 10362
rect 2786 10310 2798 10362
rect 2850 10310 2862 10362
rect 2914 10310 4078 10362
rect 4130 10310 4142 10362
rect 4194 10310 4206 10362
rect 4258 10310 4270 10362
rect 4322 10310 4334 10362
rect 4386 10310 5550 10362
rect 5602 10310 5614 10362
rect 5666 10310 5678 10362
rect 5730 10310 5742 10362
rect 5794 10310 5806 10362
rect 5858 10310 7022 10362
rect 7074 10310 7086 10362
rect 7138 10310 7150 10362
rect 7202 10310 7214 10362
rect 7266 10310 7278 10362
rect 7330 10310 7912 10362
rect 2024 10288 7912 10310
rect 6914 10208 6920 10260
rect 6972 10248 6978 10260
rect 7009 10251 7067 10257
rect 7009 10248 7021 10251
rect 6972 10220 7021 10248
rect 6972 10208 6978 10220
rect 7009 10217 7021 10220
rect 7055 10248 7067 10251
rect 7282 10248 7288 10260
rect 7055 10220 7288 10248
rect 7055 10217 7067 10220
rect 7009 10211 7067 10217
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 7374 10208 7380 10260
rect 7432 10208 7438 10260
rect 7466 10112 7472 10124
rect 6932 10084 7472 10112
rect 6932 10056 6960 10084
rect 7466 10072 7472 10084
rect 7524 10072 7530 10124
rect 6914 10004 6920 10056
rect 6972 10004 6978 10056
rect 2024 9818 8072 9840
rect 2024 9766 3342 9818
rect 3394 9766 3406 9818
rect 3458 9766 3470 9818
rect 3522 9766 3534 9818
rect 3586 9766 3598 9818
rect 3650 9766 4814 9818
rect 4866 9766 4878 9818
rect 4930 9766 4942 9818
rect 4994 9766 5006 9818
rect 5058 9766 5070 9818
rect 5122 9766 6286 9818
rect 6338 9766 6350 9818
rect 6402 9766 6414 9818
rect 6466 9766 6478 9818
rect 6530 9766 6542 9818
rect 6594 9766 7758 9818
rect 7810 9766 7822 9818
rect 7874 9766 7886 9818
rect 7938 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8072 9818
rect 2024 9744 8072 9766
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9568 7343 9571
rect 7558 9568 7564 9580
rect 7331 9540 7564 9568
rect 7331 9537 7343 9540
rect 7285 9531 7343 9537
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 7466 9392 7472 9444
rect 7524 9392 7530 9444
rect 2024 9274 7912 9296
rect 2024 9222 2606 9274
rect 2658 9222 2670 9274
rect 2722 9222 2734 9274
rect 2786 9222 2798 9274
rect 2850 9222 2862 9274
rect 2914 9222 4078 9274
rect 4130 9222 4142 9274
rect 4194 9222 4206 9274
rect 4258 9222 4270 9274
rect 4322 9222 4334 9274
rect 4386 9222 5550 9274
rect 5602 9222 5614 9274
rect 5666 9222 5678 9274
rect 5730 9222 5742 9274
rect 5794 9222 5806 9274
rect 5858 9222 7022 9274
rect 7074 9222 7086 9274
rect 7138 9222 7150 9274
rect 7202 9222 7214 9274
rect 7266 9222 7278 9274
rect 7330 9222 7912 9274
rect 2024 9200 7912 9222
rect 2024 8730 8072 8752
rect 2024 8678 3342 8730
rect 3394 8678 3406 8730
rect 3458 8678 3470 8730
rect 3522 8678 3534 8730
rect 3586 8678 3598 8730
rect 3650 8678 4814 8730
rect 4866 8678 4878 8730
rect 4930 8678 4942 8730
rect 4994 8678 5006 8730
rect 5058 8678 5070 8730
rect 5122 8678 6286 8730
rect 6338 8678 6350 8730
rect 6402 8678 6414 8730
rect 6466 8678 6478 8730
rect 6530 8678 6542 8730
rect 6594 8678 7758 8730
rect 7810 8678 7822 8730
rect 7874 8678 7886 8730
rect 7938 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8072 8730
rect 2024 8656 8072 8678
rect 2024 8186 7912 8208
rect 2024 8134 2606 8186
rect 2658 8134 2670 8186
rect 2722 8134 2734 8186
rect 2786 8134 2798 8186
rect 2850 8134 2862 8186
rect 2914 8134 4078 8186
rect 4130 8134 4142 8186
rect 4194 8134 4206 8186
rect 4258 8134 4270 8186
rect 4322 8134 4334 8186
rect 4386 8134 5550 8186
rect 5602 8134 5614 8186
rect 5666 8134 5678 8186
rect 5730 8134 5742 8186
rect 5794 8134 5806 8186
rect 5858 8134 7022 8186
rect 7074 8134 7086 8186
rect 7138 8134 7150 8186
rect 7202 8134 7214 8186
rect 7266 8134 7278 8186
rect 7330 8134 7912 8186
rect 2024 8112 7912 8134
rect 2024 7642 8072 7664
rect 2024 7590 3342 7642
rect 3394 7590 3406 7642
rect 3458 7590 3470 7642
rect 3522 7590 3534 7642
rect 3586 7590 3598 7642
rect 3650 7590 4814 7642
rect 4866 7590 4878 7642
rect 4930 7590 4942 7642
rect 4994 7590 5006 7642
rect 5058 7590 5070 7642
rect 5122 7590 6286 7642
rect 6338 7590 6350 7642
rect 6402 7590 6414 7642
rect 6466 7590 6478 7642
rect 6530 7590 6542 7642
rect 6594 7590 7758 7642
rect 7810 7590 7822 7642
rect 7874 7590 7886 7642
rect 7938 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8072 7642
rect 2024 7568 8072 7590
rect 2024 7098 7912 7120
rect 2024 7046 2606 7098
rect 2658 7046 2670 7098
rect 2722 7046 2734 7098
rect 2786 7046 2798 7098
rect 2850 7046 2862 7098
rect 2914 7046 4078 7098
rect 4130 7046 4142 7098
rect 4194 7046 4206 7098
rect 4258 7046 4270 7098
rect 4322 7046 4334 7098
rect 4386 7046 5550 7098
rect 5602 7046 5614 7098
rect 5666 7046 5678 7098
rect 5730 7046 5742 7098
rect 5794 7046 5806 7098
rect 5858 7046 7022 7098
rect 7074 7046 7086 7098
rect 7138 7046 7150 7098
rect 7202 7046 7214 7098
rect 7266 7046 7278 7098
rect 7330 7046 7912 7098
rect 2024 7024 7912 7046
rect 6914 6604 6920 6656
rect 6972 6644 6978 6656
rect 7374 6644 7380 6656
rect 6972 6616 7380 6644
rect 6972 6604 6978 6616
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 2024 6554 8072 6576
rect 2024 6502 3342 6554
rect 3394 6502 3406 6554
rect 3458 6502 3470 6554
rect 3522 6502 3534 6554
rect 3586 6502 3598 6554
rect 3650 6502 4814 6554
rect 4866 6502 4878 6554
rect 4930 6502 4942 6554
rect 4994 6502 5006 6554
rect 5058 6502 5070 6554
rect 5122 6502 6286 6554
rect 6338 6502 6350 6554
rect 6402 6502 6414 6554
rect 6466 6502 6478 6554
rect 6530 6502 6542 6554
rect 6594 6502 7758 6554
rect 7810 6502 7822 6554
rect 7874 6502 7886 6554
rect 7938 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8072 6554
rect 2024 6480 8072 6502
rect 7101 6443 7159 6449
rect 7101 6409 7113 6443
rect 7147 6409 7159 6443
rect 7101 6403 7159 6409
rect 6914 6264 6920 6316
rect 6972 6264 6978 6316
rect 7116 6304 7144 6403
rect 7285 6307 7343 6313
rect 7285 6304 7297 6307
rect 7116 6276 7297 6304
rect 7285 6273 7297 6276
rect 7331 6273 7343 6307
rect 7285 6267 7343 6273
rect 7466 6060 7472 6112
rect 7524 6060 7530 6112
rect 2024 6010 7912 6032
rect 2024 5958 2606 6010
rect 2658 5958 2670 6010
rect 2722 5958 2734 6010
rect 2786 5958 2798 6010
rect 2850 5958 2862 6010
rect 2914 5958 4078 6010
rect 4130 5958 4142 6010
rect 4194 5958 4206 6010
rect 4258 5958 4270 6010
rect 4322 5958 4334 6010
rect 4386 5958 5550 6010
rect 5602 5958 5614 6010
rect 5666 5958 5678 6010
rect 5730 5958 5742 6010
rect 5794 5958 5806 6010
rect 5858 5958 7022 6010
rect 7074 5958 7086 6010
rect 7138 5958 7150 6010
rect 7202 5958 7214 6010
rect 7266 5958 7278 6010
rect 7330 5958 7912 6010
rect 2024 5936 7912 5958
rect 6914 5856 6920 5908
rect 6972 5856 6978 5908
rect 7285 5899 7343 5905
rect 7285 5865 7297 5899
rect 7331 5896 7343 5899
rect 7374 5896 7380 5908
rect 7331 5868 7380 5896
rect 7331 5865 7343 5868
rect 7285 5859 7343 5865
rect 7374 5856 7380 5868
rect 7432 5856 7438 5908
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5692 7435 5695
rect 7558 5692 7564 5704
rect 7423 5664 7564 5692
rect 7423 5661 7435 5664
rect 7377 5655 7435 5661
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 2024 5466 8072 5488
rect 2024 5414 3342 5466
rect 3394 5414 3406 5466
rect 3458 5414 3470 5466
rect 3522 5414 3534 5466
rect 3586 5414 3598 5466
rect 3650 5414 4814 5466
rect 4866 5414 4878 5466
rect 4930 5414 4942 5466
rect 4994 5414 5006 5466
rect 5058 5414 5070 5466
rect 5122 5414 6286 5466
rect 6338 5414 6350 5466
rect 6402 5414 6414 5466
rect 6466 5414 6478 5466
rect 6530 5414 6542 5466
rect 6594 5414 7758 5466
rect 7810 5414 7822 5466
rect 7874 5414 7886 5466
rect 7938 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8072 5466
rect 2024 5392 8072 5414
rect 2024 4922 7912 4944
rect 2024 4870 2606 4922
rect 2658 4870 2670 4922
rect 2722 4870 2734 4922
rect 2786 4870 2798 4922
rect 2850 4870 2862 4922
rect 2914 4870 4078 4922
rect 4130 4870 4142 4922
rect 4194 4870 4206 4922
rect 4258 4870 4270 4922
rect 4322 4870 4334 4922
rect 4386 4870 5550 4922
rect 5602 4870 5614 4922
rect 5666 4870 5678 4922
rect 5730 4870 5742 4922
rect 5794 4870 5806 4922
rect 5858 4870 7022 4922
rect 7074 4870 7086 4922
rect 7138 4870 7150 4922
rect 7202 4870 7214 4922
rect 7266 4870 7278 4922
rect 7330 4870 7912 4922
rect 2024 4848 7912 4870
rect 2024 4378 8072 4400
rect 2024 4326 3342 4378
rect 3394 4326 3406 4378
rect 3458 4326 3470 4378
rect 3522 4326 3534 4378
rect 3586 4326 3598 4378
rect 3650 4326 4814 4378
rect 4866 4326 4878 4378
rect 4930 4326 4942 4378
rect 4994 4326 5006 4378
rect 5058 4326 5070 4378
rect 5122 4326 6286 4378
rect 6338 4326 6350 4378
rect 6402 4326 6414 4378
rect 6466 4326 6478 4378
rect 6530 4326 6542 4378
rect 6594 4326 7758 4378
rect 7810 4326 7822 4378
rect 7874 4326 7886 4378
rect 7938 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8072 4378
rect 2024 4304 8072 4326
rect 2024 3834 7912 3856
rect 2024 3782 2606 3834
rect 2658 3782 2670 3834
rect 2722 3782 2734 3834
rect 2786 3782 2798 3834
rect 2850 3782 2862 3834
rect 2914 3782 4078 3834
rect 4130 3782 4142 3834
rect 4194 3782 4206 3834
rect 4258 3782 4270 3834
rect 4322 3782 4334 3834
rect 4386 3782 5550 3834
rect 5602 3782 5614 3834
rect 5666 3782 5678 3834
rect 5730 3782 5742 3834
rect 5794 3782 5806 3834
rect 5858 3782 7022 3834
rect 7074 3782 7086 3834
rect 7138 3782 7150 3834
rect 7202 3782 7214 3834
rect 7266 3782 7278 3834
rect 7330 3782 7912 3834
rect 2024 3760 7912 3782
rect 7374 3476 7380 3528
rect 7432 3476 7438 3528
rect 7193 3451 7251 3457
rect 7193 3417 7205 3451
rect 7239 3448 7251 3451
rect 7558 3448 7564 3460
rect 7239 3420 7564 3448
rect 7239 3417 7251 3420
rect 7193 3411 7251 3417
rect 7558 3408 7564 3420
rect 7616 3408 7622 3460
rect 6638 3340 6644 3392
rect 6696 3380 6702 3392
rect 7009 3383 7067 3389
rect 7009 3380 7021 3383
rect 6696 3352 7021 3380
rect 6696 3340 6702 3352
rect 7009 3349 7021 3352
rect 7055 3349 7067 3383
rect 7009 3343 7067 3349
rect 2024 3290 8072 3312
rect 2024 3238 3342 3290
rect 3394 3238 3406 3290
rect 3458 3238 3470 3290
rect 3522 3238 3534 3290
rect 3586 3238 3598 3290
rect 3650 3238 4814 3290
rect 4866 3238 4878 3290
rect 4930 3238 4942 3290
rect 4994 3238 5006 3290
rect 5058 3238 5070 3290
rect 5122 3238 6286 3290
rect 6338 3238 6350 3290
rect 6402 3238 6414 3290
rect 6466 3238 6478 3290
rect 6530 3238 6542 3290
rect 6594 3238 7758 3290
rect 7810 3238 7822 3290
rect 7874 3238 7886 3290
rect 7938 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8072 3290
rect 2024 3216 8072 3238
rect 3145 3111 3203 3117
rect 3145 3077 3157 3111
rect 3191 3108 3203 3111
rect 7374 3108 7380 3120
rect 3191 3080 7380 3108
rect 3191 3077 3203 3080
rect 3145 3071 3203 3077
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3009 2835 3043
rect 2777 3003 2835 3009
rect 2961 3043 3019 3049
rect 2961 3009 2973 3043
rect 3007 3040 3019 3043
rect 3160 3040 3188 3071
rect 3697 3043 3755 3049
rect 3697 3040 3709 3043
rect 3007 3012 3188 3040
rect 3620 3012 3709 3040
rect 3007 3009 3019 3012
rect 2961 3003 3019 3009
rect 2792 2972 2820 3003
rect 3620 2981 3648 3012
rect 3697 3009 3709 3012
rect 3743 3009 3755 3043
rect 3697 3003 3755 3009
rect 3605 2975 3663 2981
rect 2792 2944 3556 2972
rect 3528 2913 3556 2944
rect 3605 2941 3617 2975
rect 3651 2941 3663 2975
rect 3605 2935 3663 2941
rect 5537 2975 5595 2981
rect 5537 2941 5549 2975
rect 5583 2941 5595 2975
rect 5537 2935 5595 2941
rect 3513 2907 3571 2913
rect 3513 2873 3525 2907
rect 3559 2904 3571 2907
rect 5552 2904 5580 2935
rect 5920 2913 5948 3080
rect 6089 3043 6147 3049
rect 6089 3040 6101 3043
rect 6012 3012 6101 3040
rect 6012 2981 6040 3012
rect 6089 3009 6101 3012
rect 6135 3009 6147 3043
rect 6089 3003 6147 3009
rect 6457 3043 6515 3049
rect 6457 3009 6469 3043
rect 6503 3040 6515 3043
rect 6638 3040 6644 3052
rect 6503 3012 6644 3040
rect 6503 3009 6515 3012
rect 6457 3003 6515 3009
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 6932 3049 6960 3080
rect 7374 3068 7380 3080
rect 7432 3068 7438 3120
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 7101 3043 7159 3049
rect 7101 3009 7113 3043
rect 7147 3040 7159 3043
rect 7469 3043 7527 3049
rect 7469 3040 7481 3043
rect 7147 3012 7481 3040
rect 7147 3009 7159 3012
rect 7101 3003 7159 3009
rect 7469 3009 7481 3012
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 5997 2975 6055 2981
rect 5997 2941 6009 2975
rect 6043 2941 6055 2975
rect 6733 2975 6791 2981
rect 6733 2972 6745 2975
rect 5997 2935 6055 2941
rect 6104 2944 6745 2972
rect 3559 2876 5580 2904
rect 3559 2873 3571 2876
rect 3513 2867 3571 2873
rect 2958 2796 2964 2848
rect 3016 2796 3022 2848
rect 3878 2796 3884 2848
rect 3936 2796 3942 2848
rect 5552 2836 5580 2876
rect 5905 2907 5963 2913
rect 5905 2873 5917 2907
rect 5951 2873 5963 2907
rect 5905 2867 5963 2873
rect 6104 2836 6132 2944
rect 6733 2941 6745 2944
rect 6779 2972 6791 2975
rect 7558 2972 7564 2984
rect 6779 2944 7564 2972
rect 6779 2941 6791 2944
rect 6733 2935 6791 2941
rect 7558 2932 7564 2944
rect 7616 2932 7622 2984
rect 6641 2907 6699 2913
rect 6641 2873 6653 2907
rect 6687 2904 6699 2907
rect 7374 2904 7380 2916
rect 6687 2876 7380 2904
rect 6687 2873 6699 2876
rect 6641 2867 6699 2873
rect 7374 2864 7380 2876
rect 7432 2864 7438 2916
rect 5552 2808 6132 2836
rect 6270 2796 6276 2848
rect 6328 2796 6334 2848
rect 6914 2796 6920 2848
rect 6972 2836 6978 2848
rect 7285 2839 7343 2845
rect 7285 2836 7297 2839
rect 6972 2808 7297 2836
rect 6972 2796 6978 2808
rect 7285 2805 7297 2808
rect 7331 2805 7343 2839
rect 7285 2799 7343 2805
rect 2024 2746 7912 2768
rect 2024 2694 2606 2746
rect 2658 2694 2670 2746
rect 2722 2694 2734 2746
rect 2786 2694 2798 2746
rect 2850 2694 2862 2746
rect 2914 2694 4078 2746
rect 4130 2694 4142 2746
rect 4194 2694 4206 2746
rect 4258 2694 4270 2746
rect 4322 2694 4334 2746
rect 4386 2694 5550 2746
rect 5602 2694 5614 2746
rect 5666 2694 5678 2746
rect 5730 2694 5742 2746
rect 5794 2694 5806 2746
rect 5858 2694 7022 2746
rect 7074 2694 7086 2746
rect 7138 2694 7150 2746
rect 7202 2694 7214 2746
rect 7266 2694 7278 2746
rect 7330 2694 7912 2746
rect 2024 2672 7912 2694
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2428 2743 2431
rect 2958 2428 2964 2440
rect 2731 2400 2964 2428
rect 2731 2397 2743 2400
rect 2685 2391 2743 2397
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 3878 2388 3884 2440
rect 3936 2388 3942 2440
rect 6181 2431 6239 2437
rect 6181 2397 6193 2431
rect 6227 2428 6239 2431
rect 6270 2428 6276 2440
rect 6227 2400 6276 2428
rect 6227 2397 6239 2400
rect 6181 2391 6239 2397
rect 6270 2388 6276 2400
rect 6328 2388 6334 2440
rect 6914 2388 6920 2440
rect 6972 2428 6978 2440
rect 7009 2431 7067 2437
rect 7009 2428 7021 2431
rect 6972 2400 7021 2428
rect 6972 2388 6978 2400
rect 7009 2397 7021 2400
rect 7055 2397 7067 2431
rect 7009 2391 7067 2397
rect 7285 2431 7343 2437
rect 7285 2397 7297 2431
rect 7331 2428 7343 2431
rect 7374 2428 7380 2440
rect 7331 2400 7380 2428
rect 7331 2397 7343 2400
rect 7285 2391 7343 2397
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 1210 2320 1216 2372
rect 1268 2360 1274 2372
rect 2317 2363 2375 2369
rect 2317 2360 2329 2363
rect 1268 2332 2329 2360
rect 1268 2320 1274 2332
rect 2317 2329 2329 2332
rect 2363 2329 2375 2363
rect 8662 2360 8668 2372
rect 2317 2323 2375 2329
rect 7392 2332 8668 2360
rect 3694 2252 3700 2304
rect 3752 2292 3758 2304
rect 3973 2295 4031 2301
rect 3973 2292 3985 2295
rect 3752 2264 3985 2292
rect 3752 2252 3758 2264
rect 3973 2261 3985 2264
rect 4019 2261 4031 2295
rect 3973 2255 4031 2261
rect 6178 2252 6184 2304
rect 6236 2292 6242 2304
rect 6273 2295 6331 2301
rect 6273 2292 6285 2295
rect 6236 2264 6285 2292
rect 6236 2252 6242 2264
rect 6273 2261 6285 2264
rect 6319 2261 6331 2295
rect 6273 2255 6331 2261
rect 6917 2295 6975 2301
rect 6917 2261 6929 2295
rect 6963 2292 6975 2295
rect 7392 2292 7420 2332
rect 8662 2320 8668 2332
rect 8720 2320 8726 2372
rect 6963 2264 7420 2292
rect 7469 2295 7527 2301
rect 6963 2261 6975 2264
rect 6917 2255 6975 2261
rect 7469 2261 7481 2295
rect 7515 2292 7527 2295
rect 8202 2292 8208 2304
rect 7515 2264 8208 2292
rect 7515 2261 7527 2264
rect 7469 2255 7527 2261
rect 8202 2252 8208 2264
rect 8260 2252 8266 2304
rect 2024 2202 8072 2224
rect 2024 2150 3342 2202
rect 3394 2150 3406 2202
rect 3458 2150 3470 2202
rect 3522 2150 3534 2202
rect 3586 2150 3598 2202
rect 3650 2150 4814 2202
rect 4866 2150 4878 2202
rect 4930 2150 4942 2202
rect 4994 2150 5006 2202
rect 5058 2150 5070 2202
rect 5122 2150 6286 2202
rect 6338 2150 6350 2202
rect 6402 2150 6414 2202
rect 6466 2150 6478 2202
rect 6530 2150 6542 2202
rect 6594 2150 7758 2202
rect 7810 2150 7822 2202
rect 7874 2150 7886 2202
rect 7938 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8072 2202
rect 2024 2128 8072 2150
<< via1 >>
rect 2606 13574 2658 13626
rect 2670 13574 2722 13626
rect 2734 13574 2786 13626
rect 2798 13574 2850 13626
rect 2862 13574 2914 13626
rect 4078 13574 4130 13626
rect 4142 13574 4194 13626
rect 4206 13574 4258 13626
rect 4270 13574 4322 13626
rect 4334 13574 4386 13626
rect 5550 13574 5602 13626
rect 5614 13574 5666 13626
rect 5678 13574 5730 13626
rect 5742 13574 5794 13626
rect 5806 13574 5858 13626
rect 7022 13574 7074 13626
rect 7086 13574 7138 13626
rect 7150 13574 7202 13626
rect 7214 13574 7266 13626
rect 7278 13574 7330 13626
rect 8300 13404 8352 13456
rect 2504 13268 2556 13320
rect 7472 13311 7524 13320
rect 7472 13277 7481 13311
rect 7481 13277 7515 13311
rect 7515 13277 7524 13311
rect 7472 13268 7524 13277
rect 6920 13200 6972 13252
rect 7288 13200 7340 13252
rect 7472 13132 7524 13184
rect 3342 13030 3394 13082
rect 3406 13030 3458 13082
rect 3470 13030 3522 13082
rect 3534 13030 3586 13082
rect 3598 13030 3650 13082
rect 4814 13030 4866 13082
rect 4878 13030 4930 13082
rect 4942 13030 4994 13082
rect 5006 13030 5058 13082
rect 5070 13030 5122 13082
rect 6286 13030 6338 13082
rect 6350 13030 6402 13082
rect 6414 13030 6466 13082
rect 6478 13030 6530 13082
rect 6542 13030 6594 13082
rect 7758 13030 7810 13082
rect 7822 13030 7874 13082
rect 7886 13030 7938 13082
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 7288 12971 7340 12980
rect 7288 12937 7297 12971
rect 7297 12937 7331 12971
rect 7331 12937 7340 12971
rect 7288 12928 7340 12937
rect 6920 12792 6972 12844
rect 7472 12835 7524 12844
rect 7472 12801 7481 12835
rect 7481 12801 7515 12835
rect 7515 12801 7524 12835
rect 7472 12792 7524 12801
rect 2606 12486 2658 12538
rect 2670 12486 2722 12538
rect 2734 12486 2786 12538
rect 2798 12486 2850 12538
rect 2862 12486 2914 12538
rect 4078 12486 4130 12538
rect 4142 12486 4194 12538
rect 4206 12486 4258 12538
rect 4270 12486 4322 12538
rect 4334 12486 4386 12538
rect 5550 12486 5602 12538
rect 5614 12486 5666 12538
rect 5678 12486 5730 12538
rect 5742 12486 5794 12538
rect 5806 12486 5858 12538
rect 7022 12486 7074 12538
rect 7086 12486 7138 12538
rect 7150 12486 7202 12538
rect 7214 12486 7266 12538
rect 7278 12486 7330 12538
rect 3342 11942 3394 11994
rect 3406 11942 3458 11994
rect 3470 11942 3522 11994
rect 3534 11942 3586 11994
rect 3598 11942 3650 11994
rect 4814 11942 4866 11994
rect 4878 11942 4930 11994
rect 4942 11942 4994 11994
rect 5006 11942 5058 11994
rect 5070 11942 5122 11994
rect 6286 11942 6338 11994
rect 6350 11942 6402 11994
rect 6414 11942 6466 11994
rect 6478 11942 6530 11994
rect 6542 11942 6594 11994
rect 7758 11942 7810 11994
rect 7822 11942 7874 11994
rect 7886 11942 7938 11994
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 2606 11398 2658 11450
rect 2670 11398 2722 11450
rect 2734 11398 2786 11450
rect 2798 11398 2850 11450
rect 2862 11398 2914 11450
rect 4078 11398 4130 11450
rect 4142 11398 4194 11450
rect 4206 11398 4258 11450
rect 4270 11398 4322 11450
rect 4334 11398 4386 11450
rect 5550 11398 5602 11450
rect 5614 11398 5666 11450
rect 5678 11398 5730 11450
rect 5742 11398 5794 11450
rect 5806 11398 5858 11450
rect 7022 11398 7074 11450
rect 7086 11398 7138 11450
rect 7150 11398 7202 11450
rect 7214 11398 7266 11450
rect 7278 11398 7330 11450
rect 3342 10854 3394 10906
rect 3406 10854 3458 10906
rect 3470 10854 3522 10906
rect 3534 10854 3586 10906
rect 3598 10854 3650 10906
rect 4814 10854 4866 10906
rect 4878 10854 4930 10906
rect 4942 10854 4994 10906
rect 5006 10854 5058 10906
rect 5070 10854 5122 10906
rect 6286 10854 6338 10906
rect 6350 10854 6402 10906
rect 6414 10854 6466 10906
rect 6478 10854 6530 10906
rect 6542 10854 6594 10906
rect 7758 10854 7810 10906
rect 7822 10854 7874 10906
rect 7886 10854 7938 10906
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 7380 10616 7432 10668
rect 7564 10412 7616 10464
rect 2606 10310 2658 10362
rect 2670 10310 2722 10362
rect 2734 10310 2786 10362
rect 2798 10310 2850 10362
rect 2862 10310 2914 10362
rect 4078 10310 4130 10362
rect 4142 10310 4194 10362
rect 4206 10310 4258 10362
rect 4270 10310 4322 10362
rect 4334 10310 4386 10362
rect 5550 10310 5602 10362
rect 5614 10310 5666 10362
rect 5678 10310 5730 10362
rect 5742 10310 5794 10362
rect 5806 10310 5858 10362
rect 7022 10310 7074 10362
rect 7086 10310 7138 10362
rect 7150 10310 7202 10362
rect 7214 10310 7266 10362
rect 7278 10310 7330 10362
rect 6920 10208 6972 10260
rect 7288 10208 7340 10260
rect 7380 10251 7432 10260
rect 7380 10217 7389 10251
rect 7389 10217 7423 10251
rect 7423 10217 7432 10251
rect 7380 10208 7432 10217
rect 7472 10072 7524 10124
rect 6920 10047 6972 10056
rect 6920 10013 6929 10047
rect 6929 10013 6963 10047
rect 6963 10013 6972 10047
rect 6920 10004 6972 10013
rect 3342 9766 3394 9818
rect 3406 9766 3458 9818
rect 3470 9766 3522 9818
rect 3534 9766 3586 9818
rect 3598 9766 3650 9818
rect 4814 9766 4866 9818
rect 4878 9766 4930 9818
rect 4942 9766 4994 9818
rect 5006 9766 5058 9818
rect 5070 9766 5122 9818
rect 6286 9766 6338 9818
rect 6350 9766 6402 9818
rect 6414 9766 6466 9818
rect 6478 9766 6530 9818
rect 6542 9766 6594 9818
rect 7758 9766 7810 9818
rect 7822 9766 7874 9818
rect 7886 9766 7938 9818
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 7564 9528 7616 9580
rect 7472 9435 7524 9444
rect 7472 9401 7481 9435
rect 7481 9401 7515 9435
rect 7515 9401 7524 9435
rect 7472 9392 7524 9401
rect 2606 9222 2658 9274
rect 2670 9222 2722 9274
rect 2734 9222 2786 9274
rect 2798 9222 2850 9274
rect 2862 9222 2914 9274
rect 4078 9222 4130 9274
rect 4142 9222 4194 9274
rect 4206 9222 4258 9274
rect 4270 9222 4322 9274
rect 4334 9222 4386 9274
rect 5550 9222 5602 9274
rect 5614 9222 5666 9274
rect 5678 9222 5730 9274
rect 5742 9222 5794 9274
rect 5806 9222 5858 9274
rect 7022 9222 7074 9274
rect 7086 9222 7138 9274
rect 7150 9222 7202 9274
rect 7214 9222 7266 9274
rect 7278 9222 7330 9274
rect 3342 8678 3394 8730
rect 3406 8678 3458 8730
rect 3470 8678 3522 8730
rect 3534 8678 3586 8730
rect 3598 8678 3650 8730
rect 4814 8678 4866 8730
rect 4878 8678 4930 8730
rect 4942 8678 4994 8730
rect 5006 8678 5058 8730
rect 5070 8678 5122 8730
rect 6286 8678 6338 8730
rect 6350 8678 6402 8730
rect 6414 8678 6466 8730
rect 6478 8678 6530 8730
rect 6542 8678 6594 8730
rect 7758 8678 7810 8730
rect 7822 8678 7874 8730
rect 7886 8678 7938 8730
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 2606 8134 2658 8186
rect 2670 8134 2722 8186
rect 2734 8134 2786 8186
rect 2798 8134 2850 8186
rect 2862 8134 2914 8186
rect 4078 8134 4130 8186
rect 4142 8134 4194 8186
rect 4206 8134 4258 8186
rect 4270 8134 4322 8186
rect 4334 8134 4386 8186
rect 5550 8134 5602 8186
rect 5614 8134 5666 8186
rect 5678 8134 5730 8186
rect 5742 8134 5794 8186
rect 5806 8134 5858 8186
rect 7022 8134 7074 8186
rect 7086 8134 7138 8186
rect 7150 8134 7202 8186
rect 7214 8134 7266 8186
rect 7278 8134 7330 8186
rect 3342 7590 3394 7642
rect 3406 7590 3458 7642
rect 3470 7590 3522 7642
rect 3534 7590 3586 7642
rect 3598 7590 3650 7642
rect 4814 7590 4866 7642
rect 4878 7590 4930 7642
rect 4942 7590 4994 7642
rect 5006 7590 5058 7642
rect 5070 7590 5122 7642
rect 6286 7590 6338 7642
rect 6350 7590 6402 7642
rect 6414 7590 6466 7642
rect 6478 7590 6530 7642
rect 6542 7590 6594 7642
rect 7758 7590 7810 7642
rect 7822 7590 7874 7642
rect 7886 7590 7938 7642
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 2606 7046 2658 7098
rect 2670 7046 2722 7098
rect 2734 7046 2786 7098
rect 2798 7046 2850 7098
rect 2862 7046 2914 7098
rect 4078 7046 4130 7098
rect 4142 7046 4194 7098
rect 4206 7046 4258 7098
rect 4270 7046 4322 7098
rect 4334 7046 4386 7098
rect 5550 7046 5602 7098
rect 5614 7046 5666 7098
rect 5678 7046 5730 7098
rect 5742 7046 5794 7098
rect 5806 7046 5858 7098
rect 7022 7046 7074 7098
rect 7086 7046 7138 7098
rect 7150 7046 7202 7098
rect 7214 7046 7266 7098
rect 7278 7046 7330 7098
rect 6920 6604 6972 6656
rect 7380 6604 7432 6656
rect 3342 6502 3394 6554
rect 3406 6502 3458 6554
rect 3470 6502 3522 6554
rect 3534 6502 3586 6554
rect 3598 6502 3650 6554
rect 4814 6502 4866 6554
rect 4878 6502 4930 6554
rect 4942 6502 4994 6554
rect 5006 6502 5058 6554
rect 5070 6502 5122 6554
rect 6286 6502 6338 6554
rect 6350 6502 6402 6554
rect 6414 6502 6466 6554
rect 6478 6502 6530 6554
rect 6542 6502 6594 6554
rect 7758 6502 7810 6554
rect 7822 6502 7874 6554
rect 7886 6502 7938 6554
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 6920 6307 6972 6316
rect 6920 6273 6929 6307
rect 6929 6273 6963 6307
rect 6963 6273 6972 6307
rect 6920 6264 6972 6273
rect 7472 6103 7524 6112
rect 7472 6069 7481 6103
rect 7481 6069 7515 6103
rect 7515 6069 7524 6103
rect 7472 6060 7524 6069
rect 2606 5958 2658 6010
rect 2670 5958 2722 6010
rect 2734 5958 2786 6010
rect 2798 5958 2850 6010
rect 2862 5958 2914 6010
rect 4078 5958 4130 6010
rect 4142 5958 4194 6010
rect 4206 5958 4258 6010
rect 4270 5958 4322 6010
rect 4334 5958 4386 6010
rect 5550 5958 5602 6010
rect 5614 5958 5666 6010
rect 5678 5958 5730 6010
rect 5742 5958 5794 6010
rect 5806 5958 5858 6010
rect 7022 5958 7074 6010
rect 7086 5958 7138 6010
rect 7150 5958 7202 6010
rect 7214 5958 7266 6010
rect 7278 5958 7330 6010
rect 6920 5899 6972 5908
rect 6920 5865 6929 5899
rect 6929 5865 6963 5899
rect 6963 5865 6972 5899
rect 6920 5856 6972 5865
rect 7380 5856 7432 5908
rect 7564 5652 7616 5704
rect 3342 5414 3394 5466
rect 3406 5414 3458 5466
rect 3470 5414 3522 5466
rect 3534 5414 3586 5466
rect 3598 5414 3650 5466
rect 4814 5414 4866 5466
rect 4878 5414 4930 5466
rect 4942 5414 4994 5466
rect 5006 5414 5058 5466
rect 5070 5414 5122 5466
rect 6286 5414 6338 5466
rect 6350 5414 6402 5466
rect 6414 5414 6466 5466
rect 6478 5414 6530 5466
rect 6542 5414 6594 5466
rect 7758 5414 7810 5466
rect 7822 5414 7874 5466
rect 7886 5414 7938 5466
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 2606 4870 2658 4922
rect 2670 4870 2722 4922
rect 2734 4870 2786 4922
rect 2798 4870 2850 4922
rect 2862 4870 2914 4922
rect 4078 4870 4130 4922
rect 4142 4870 4194 4922
rect 4206 4870 4258 4922
rect 4270 4870 4322 4922
rect 4334 4870 4386 4922
rect 5550 4870 5602 4922
rect 5614 4870 5666 4922
rect 5678 4870 5730 4922
rect 5742 4870 5794 4922
rect 5806 4870 5858 4922
rect 7022 4870 7074 4922
rect 7086 4870 7138 4922
rect 7150 4870 7202 4922
rect 7214 4870 7266 4922
rect 7278 4870 7330 4922
rect 3342 4326 3394 4378
rect 3406 4326 3458 4378
rect 3470 4326 3522 4378
rect 3534 4326 3586 4378
rect 3598 4326 3650 4378
rect 4814 4326 4866 4378
rect 4878 4326 4930 4378
rect 4942 4326 4994 4378
rect 5006 4326 5058 4378
rect 5070 4326 5122 4378
rect 6286 4326 6338 4378
rect 6350 4326 6402 4378
rect 6414 4326 6466 4378
rect 6478 4326 6530 4378
rect 6542 4326 6594 4378
rect 7758 4326 7810 4378
rect 7822 4326 7874 4378
rect 7886 4326 7938 4378
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 2606 3782 2658 3834
rect 2670 3782 2722 3834
rect 2734 3782 2786 3834
rect 2798 3782 2850 3834
rect 2862 3782 2914 3834
rect 4078 3782 4130 3834
rect 4142 3782 4194 3834
rect 4206 3782 4258 3834
rect 4270 3782 4322 3834
rect 4334 3782 4386 3834
rect 5550 3782 5602 3834
rect 5614 3782 5666 3834
rect 5678 3782 5730 3834
rect 5742 3782 5794 3834
rect 5806 3782 5858 3834
rect 7022 3782 7074 3834
rect 7086 3782 7138 3834
rect 7150 3782 7202 3834
rect 7214 3782 7266 3834
rect 7278 3782 7330 3834
rect 7380 3519 7432 3528
rect 7380 3485 7389 3519
rect 7389 3485 7423 3519
rect 7423 3485 7432 3519
rect 7380 3476 7432 3485
rect 7564 3408 7616 3460
rect 6644 3340 6696 3392
rect 3342 3238 3394 3290
rect 3406 3238 3458 3290
rect 3470 3238 3522 3290
rect 3534 3238 3586 3290
rect 3598 3238 3650 3290
rect 4814 3238 4866 3290
rect 4878 3238 4930 3290
rect 4942 3238 4994 3290
rect 5006 3238 5058 3290
rect 5070 3238 5122 3290
rect 6286 3238 6338 3290
rect 6350 3238 6402 3290
rect 6414 3238 6466 3290
rect 6478 3238 6530 3290
rect 6542 3238 6594 3290
rect 7758 3238 7810 3290
rect 7822 3238 7874 3290
rect 7886 3238 7938 3290
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 6644 3000 6696 3052
rect 7380 3068 7432 3120
rect 2964 2839 3016 2848
rect 2964 2805 2973 2839
rect 2973 2805 3007 2839
rect 3007 2805 3016 2839
rect 2964 2796 3016 2805
rect 3884 2839 3936 2848
rect 3884 2805 3893 2839
rect 3893 2805 3927 2839
rect 3927 2805 3936 2839
rect 3884 2796 3936 2805
rect 7564 2932 7616 2984
rect 7380 2864 7432 2916
rect 6276 2839 6328 2848
rect 6276 2805 6285 2839
rect 6285 2805 6319 2839
rect 6319 2805 6328 2839
rect 6276 2796 6328 2805
rect 6920 2796 6972 2848
rect 2606 2694 2658 2746
rect 2670 2694 2722 2746
rect 2734 2694 2786 2746
rect 2798 2694 2850 2746
rect 2862 2694 2914 2746
rect 4078 2694 4130 2746
rect 4142 2694 4194 2746
rect 4206 2694 4258 2746
rect 4270 2694 4322 2746
rect 4334 2694 4386 2746
rect 5550 2694 5602 2746
rect 5614 2694 5666 2746
rect 5678 2694 5730 2746
rect 5742 2694 5794 2746
rect 5806 2694 5858 2746
rect 7022 2694 7074 2746
rect 7086 2694 7138 2746
rect 7150 2694 7202 2746
rect 7214 2694 7266 2746
rect 7278 2694 7330 2746
rect 2964 2388 3016 2440
rect 3884 2431 3936 2440
rect 3884 2397 3893 2431
rect 3893 2397 3927 2431
rect 3927 2397 3936 2431
rect 3884 2388 3936 2397
rect 6276 2388 6328 2440
rect 6920 2388 6972 2440
rect 7380 2388 7432 2440
rect 1216 2320 1268 2372
rect 3700 2252 3752 2304
rect 6184 2252 6236 2304
rect 8668 2320 8720 2372
rect 8208 2252 8260 2304
rect 3342 2150 3394 2202
rect 3406 2150 3458 2202
rect 3470 2150 3522 2202
rect 3534 2150 3586 2202
rect 3598 2150 3650 2202
rect 4814 2150 4866 2202
rect 4878 2150 4930 2202
rect 4942 2150 4994 2202
rect 5006 2150 5058 2202
rect 5070 2150 5122 2202
rect 6286 2150 6338 2202
rect 6350 2150 6402 2202
rect 6414 2150 6466 2202
rect 6478 2150 6530 2202
rect 6542 2150 6594 2202
rect 7758 2150 7810 2202
rect 7822 2150 7874 2202
rect 7886 2150 7938 2202
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
<< metal2 >>
rect 2502 15600 2558 16000
rect 7470 15600 7526 16000
rect 2516 13326 2544 15600
rect 2606 13628 2914 13637
rect 2606 13626 2612 13628
rect 2668 13626 2692 13628
rect 2748 13626 2772 13628
rect 2828 13626 2852 13628
rect 2908 13626 2914 13628
rect 2668 13574 2670 13626
rect 2850 13574 2852 13626
rect 2606 13572 2612 13574
rect 2668 13572 2692 13574
rect 2748 13572 2772 13574
rect 2828 13572 2852 13574
rect 2908 13572 2914 13574
rect 2606 13563 2914 13572
rect 4078 13628 4386 13637
rect 4078 13626 4084 13628
rect 4140 13626 4164 13628
rect 4220 13626 4244 13628
rect 4300 13626 4324 13628
rect 4380 13626 4386 13628
rect 4140 13574 4142 13626
rect 4322 13574 4324 13626
rect 4078 13572 4084 13574
rect 4140 13572 4164 13574
rect 4220 13572 4244 13574
rect 4300 13572 4324 13574
rect 4380 13572 4386 13574
rect 4078 13563 4386 13572
rect 5550 13628 5858 13637
rect 5550 13626 5556 13628
rect 5612 13626 5636 13628
rect 5692 13626 5716 13628
rect 5772 13626 5796 13628
rect 5852 13626 5858 13628
rect 5612 13574 5614 13626
rect 5794 13574 5796 13626
rect 5550 13572 5556 13574
rect 5612 13572 5636 13574
rect 5692 13572 5716 13574
rect 5772 13572 5796 13574
rect 5852 13572 5858 13574
rect 5550 13563 5858 13572
rect 7022 13628 7330 13637
rect 7022 13626 7028 13628
rect 7084 13626 7108 13628
rect 7164 13626 7188 13628
rect 7244 13626 7268 13628
rect 7324 13626 7330 13628
rect 7084 13574 7086 13626
rect 7266 13574 7268 13626
rect 7022 13572 7028 13574
rect 7084 13572 7108 13574
rect 7164 13572 7188 13574
rect 7244 13572 7268 13574
rect 7324 13572 7330 13574
rect 7022 13563 7330 13572
rect 7484 13326 7512 15600
rect 8298 13696 8354 13705
rect 8298 13631 8354 13640
rect 8312 13462 8340 13631
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 3342 13084 3650 13093
rect 3342 13082 3348 13084
rect 3404 13082 3428 13084
rect 3484 13082 3508 13084
rect 3564 13082 3588 13084
rect 3644 13082 3650 13084
rect 3404 13030 3406 13082
rect 3586 13030 3588 13082
rect 3342 13028 3348 13030
rect 3404 13028 3428 13030
rect 3484 13028 3508 13030
rect 3564 13028 3588 13030
rect 3644 13028 3650 13030
rect 3342 13019 3650 13028
rect 4814 13084 5122 13093
rect 4814 13082 4820 13084
rect 4876 13082 4900 13084
rect 4956 13082 4980 13084
rect 5036 13082 5060 13084
rect 5116 13082 5122 13084
rect 4876 13030 4878 13082
rect 5058 13030 5060 13082
rect 4814 13028 4820 13030
rect 4876 13028 4900 13030
rect 4956 13028 4980 13030
rect 5036 13028 5060 13030
rect 5116 13028 5122 13030
rect 4814 13019 5122 13028
rect 6286 13084 6594 13093
rect 6286 13082 6292 13084
rect 6348 13082 6372 13084
rect 6428 13082 6452 13084
rect 6508 13082 6532 13084
rect 6588 13082 6594 13084
rect 6348 13030 6350 13082
rect 6530 13030 6532 13082
rect 6286 13028 6292 13030
rect 6348 13028 6372 13030
rect 6428 13028 6452 13030
rect 6508 13028 6532 13030
rect 6588 13028 6594 13030
rect 6286 13019 6594 13028
rect 6932 12850 6960 13194
rect 7300 12986 7328 13194
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7484 12850 7512 13126
rect 7758 13084 8066 13093
rect 7758 13082 7764 13084
rect 7820 13082 7844 13084
rect 7900 13082 7924 13084
rect 7980 13082 8004 13084
rect 8060 13082 8066 13084
rect 7820 13030 7822 13082
rect 8002 13030 8004 13082
rect 7758 13028 7764 13030
rect 7820 13028 7844 13030
rect 7900 13028 7924 13030
rect 7980 13028 8004 13030
rect 8060 13028 8066 13030
rect 7758 13019 8066 13028
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 2606 12540 2914 12549
rect 2606 12538 2612 12540
rect 2668 12538 2692 12540
rect 2748 12538 2772 12540
rect 2828 12538 2852 12540
rect 2908 12538 2914 12540
rect 2668 12486 2670 12538
rect 2850 12486 2852 12538
rect 2606 12484 2612 12486
rect 2668 12484 2692 12486
rect 2748 12484 2772 12486
rect 2828 12484 2852 12486
rect 2908 12484 2914 12486
rect 2606 12475 2914 12484
rect 4078 12540 4386 12549
rect 4078 12538 4084 12540
rect 4140 12538 4164 12540
rect 4220 12538 4244 12540
rect 4300 12538 4324 12540
rect 4380 12538 4386 12540
rect 4140 12486 4142 12538
rect 4322 12486 4324 12538
rect 4078 12484 4084 12486
rect 4140 12484 4164 12486
rect 4220 12484 4244 12486
rect 4300 12484 4324 12486
rect 4380 12484 4386 12486
rect 4078 12475 4386 12484
rect 5550 12540 5858 12549
rect 5550 12538 5556 12540
rect 5612 12538 5636 12540
rect 5692 12538 5716 12540
rect 5772 12538 5796 12540
rect 5852 12538 5858 12540
rect 5612 12486 5614 12538
rect 5794 12486 5796 12538
rect 5550 12484 5556 12486
rect 5612 12484 5636 12486
rect 5692 12484 5716 12486
rect 5772 12484 5796 12486
rect 5852 12484 5858 12486
rect 5550 12475 5858 12484
rect 3342 11996 3650 12005
rect 3342 11994 3348 11996
rect 3404 11994 3428 11996
rect 3484 11994 3508 11996
rect 3564 11994 3588 11996
rect 3644 11994 3650 11996
rect 3404 11942 3406 11994
rect 3586 11942 3588 11994
rect 3342 11940 3348 11942
rect 3404 11940 3428 11942
rect 3484 11940 3508 11942
rect 3564 11940 3588 11942
rect 3644 11940 3650 11942
rect 3342 11931 3650 11940
rect 4814 11996 5122 12005
rect 4814 11994 4820 11996
rect 4876 11994 4900 11996
rect 4956 11994 4980 11996
rect 5036 11994 5060 11996
rect 5116 11994 5122 11996
rect 4876 11942 4878 11994
rect 5058 11942 5060 11994
rect 4814 11940 4820 11942
rect 4876 11940 4900 11942
rect 4956 11940 4980 11942
rect 5036 11940 5060 11942
rect 5116 11940 5122 11942
rect 4814 11931 5122 11940
rect 6286 11996 6594 12005
rect 6286 11994 6292 11996
rect 6348 11994 6372 11996
rect 6428 11994 6452 11996
rect 6508 11994 6532 11996
rect 6588 11994 6594 11996
rect 6348 11942 6350 11994
rect 6530 11942 6532 11994
rect 6286 11940 6292 11942
rect 6348 11940 6372 11942
rect 6428 11940 6452 11942
rect 6508 11940 6532 11942
rect 6588 11940 6594 11942
rect 6286 11931 6594 11940
rect 2606 11452 2914 11461
rect 2606 11450 2612 11452
rect 2668 11450 2692 11452
rect 2748 11450 2772 11452
rect 2828 11450 2852 11452
rect 2908 11450 2914 11452
rect 2668 11398 2670 11450
rect 2850 11398 2852 11450
rect 2606 11396 2612 11398
rect 2668 11396 2692 11398
rect 2748 11396 2772 11398
rect 2828 11396 2852 11398
rect 2908 11396 2914 11398
rect 2606 11387 2914 11396
rect 4078 11452 4386 11461
rect 4078 11450 4084 11452
rect 4140 11450 4164 11452
rect 4220 11450 4244 11452
rect 4300 11450 4324 11452
rect 4380 11450 4386 11452
rect 4140 11398 4142 11450
rect 4322 11398 4324 11450
rect 4078 11396 4084 11398
rect 4140 11396 4164 11398
rect 4220 11396 4244 11398
rect 4300 11396 4324 11398
rect 4380 11396 4386 11398
rect 4078 11387 4386 11396
rect 5550 11452 5858 11461
rect 5550 11450 5556 11452
rect 5612 11450 5636 11452
rect 5692 11450 5716 11452
rect 5772 11450 5796 11452
rect 5852 11450 5858 11452
rect 5612 11398 5614 11450
rect 5794 11398 5796 11450
rect 5550 11396 5556 11398
rect 5612 11396 5636 11398
rect 5692 11396 5716 11398
rect 5772 11396 5796 11398
rect 5852 11396 5858 11398
rect 5550 11387 5858 11396
rect 3342 10908 3650 10917
rect 3342 10906 3348 10908
rect 3404 10906 3428 10908
rect 3484 10906 3508 10908
rect 3564 10906 3588 10908
rect 3644 10906 3650 10908
rect 3404 10854 3406 10906
rect 3586 10854 3588 10906
rect 3342 10852 3348 10854
rect 3404 10852 3428 10854
rect 3484 10852 3508 10854
rect 3564 10852 3588 10854
rect 3644 10852 3650 10854
rect 3342 10843 3650 10852
rect 4814 10908 5122 10917
rect 4814 10906 4820 10908
rect 4876 10906 4900 10908
rect 4956 10906 4980 10908
rect 5036 10906 5060 10908
rect 5116 10906 5122 10908
rect 4876 10854 4878 10906
rect 5058 10854 5060 10906
rect 4814 10852 4820 10854
rect 4876 10852 4900 10854
rect 4956 10852 4980 10854
rect 5036 10852 5060 10854
rect 5116 10852 5122 10854
rect 4814 10843 5122 10852
rect 6286 10908 6594 10917
rect 6286 10906 6292 10908
rect 6348 10906 6372 10908
rect 6428 10906 6452 10908
rect 6508 10906 6532 10908
rect 6588 10906 6594 10908
rect 6348 10854 6350 10906
rect 6530 10854 6532 10906
rect 6286 10852 6292 10854
rect 6348 10852 6372 10854
rect 6428 10852 6452 10854
rect 6508 10852 6532 10854
rect 6588 10852 6594 10854
rect 6286 10843 6594 10852
rect 2606 10364 2914 10373
rect 2606 10362 2612 10364
rect 2668 10362 2692 10364
rect 2748 10362 2772 10364
rect 2828 10362 2852 10364
rect 2908 10362 2914 10364
rect 2668 10310 2670 10362
rect 2850 10310 2852 10362
rect 2606 10308 2612 10310
rect 2668 10308 2692 10310
rect 2748 10308 2772 10310
rect 2828 10308 2852 10310
rect 2908 10308 2914 10310
rect 2606 10299 2914 10308
rect 4078 10364 4386 10373
rect 4078 10362 4084 10364
rect 4140 10362 4164 10364
rect 4220 10362 4244 10364
rect 4300 10362 4324 10364
rect 4380 10362 4386 10364
rect 4140 10310 4142 10362
rect 4322 10310 4324 10362
rect 4078 10308 4084 10310
rect 4140 10308 4164 10310
rect 4220 10308 4244 10310
rect 4300 10308 4324 10310
rect 4380 10308 4386 10310
rect 4078 10299 4386 10308
rect 5550 10364 5858 10373
rect 5550 10362 5556 10364
rect 5612 10362 5636 10364
rect 5692 10362 5716 10364
rect 5772 10362 5796 10364
rect 5852 10362 5858 10364
rect 5612 10310 5614 10362
rect 5794 10310 5796 10362
rect 5550 10308 5556 10310
rect 5612 10308 5636 10310
rect 5692 10308 5716 10310
rect 5772 10308 5796 10310
rect 5852 10308 5858 10310
rect 5550 10299 5858 10308
rect 6932 10266 6960 12786
rect 7022 12540 7330 12549
rect 7022 12538 7028 12540
rect 7084 12538 7108 12540
rect 7164 12538 7188 12540
rect 7244 12538 7268 12540
rect 7324 12538 7330 12540
rect 7084 12486 7086 12538
rect 7266 12486 7268 12538
rect 7022 12484 7028 12486
rect 7084 12484 7108 12486
rect 7164 12484 7188 12486
rect 7244 12484 7268 12486
rect 7324 12484 7330 12486
rect 7022 12475 7330 12484
rect 7022 11452 7330 11461
rect 7022 11450 7028 11452
rect 7084 11450 7108 11452
rect 7164 11450 7188 11452
rect 7244 11450 7268 11452
rect 7324 11450 7330 11452
rect 7084 11398 7086 11450
rect 7266 11398 7268 11450
rect 7022 11396 7028 11398
rect 7084 11396 7108 11398
rect 7164 11396 7188 11398
rect 7244 11396 7268 11398
rect 7324 11396 7330 11398
rect 7022 11387 7330 11396
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7022 10364 7330 10373
rect 7022 10362 7028 10364
rect 7084 10362 7108 10364
rect 7164 10362 7188 10364
rect 7244 10362 7268 10364
rect 7324 10362 7330 10364
rect 7084 10310 7086 10362
rect 7266 10310 7268 10362
rect 7022 10308 7028 10310
rect 7084 10308 7108 10310
rect 7164 10308 7188 10310
rect 7244 10308 7268 10310
rect 7324 10308 7330 10310
rect 7022 10299 7330 10308
rect 7392 10266 7420 10610
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 3342 9820 3650 9829
rect 3342 9818 3348 9820
rect 3404 9818 3428 9820
rect 3484 9818 3508 9820
rect 3564 9818 3588 9820
rect 3644 9818 3650 9820
rect 3404 9766 3406 9818
rect 3586 9766 3588 9818
rect 3342 9764 3348 9766
rect 3404 9764 3428 9766
rect 3484 9764 3508 9766
rect 3564 9764 3588 9766
rect 3644 9764 3650 9766
rect 3342 9755 3650 9764
rect 4814 9820 5122 9829
rect 4814 9818 4820 9820
rect 4876 9818 4900 9820
rect 4956 9818 4980 9820
rect 5036 9818 5060 9820
rect 5116 9818 5122 9820
rect 4876 9766 4878 9818
rect 5058 9766 5060 9818
rect 4814 9764 4820 9766
rect 4876 9764 4900 9766
rect 4956 9764 4980 9766
rect 5036 9764 5060 9766
rect 5116 9764 5122 9766
rect 4814 9755 5122 9764
rect 6286 9820 6594 9829
rect 6286 9818 6292 9820
rect 6348 9818 6372 9820
rect 6428 9818 6452 9820
rect 6508 9818 6532 9820
rect 6588 9818 6594 9820
rect 6348 9766 6350 9818
rect 6530 9766 6532 9818
rect 6286 9764 6292 9766
rect 6348 9764 6372 9766
rect 6428 9764 6452 9766
rect 6508 9764 6532 9766
rect 6588 9764 6594 9766
rect 6286 9755 6594 9764
rect 2606 9276 2914 9285
rect 2606 9274 2612 9276
rect 2668 9274 2692 9276
rect 2748 9274 2772 9276
rect 2828 9274 2852 9276
rect 2908 9274 2914 9276
rect 2668 9222 2670 9274
rect 2850 9222 2852 9274
rect 2606 9220 2612 9222
rect 2668 9220 2692 9222
rect 2748 9220 2772 9222
rect 2828 9220 2852 9222
rect 2908 9220 2914 9222
rect 2606 9211 2914 9220
rect 4078 9276 4386 9285
rect 4078 9274 4084 9276
rect 4140 9274 4164 9276
rect 4220 9274 4244 9276
rect 4300 9274 4324 9276
rect 4380 9274 4386 9276
rect 4140 9222 4142 9274
rect 4322 9222 4324 9274
rect 4078 9220 4084 9222
rect 4140 9220 4164 9222
rect 4220 9220 4244 9222
rect 4300 9220 4324 9222
rect 4380 9220 4386 9222
rect 4078 9211 4386 9220
rect 5550 9276 5858 9285
rect 5550 9274 5556 9276
rect 5612 9274 5636 9276
rect 5692 9274 5716 9276
rect 5772 9274 5796 9276
rect 5852 9274 5858 9276
rect 5612 9222 5614 9274
rect 5794 9222 5796 9274
rect 5550 9220 5556 9222
rect 5612 9220 5636 9222
rect 5692 9220 5716 9222
rect 5772 9220 5796 9222
rect 5852 9220 5858 9222
rect 5550 9211 5858 9220
rect 3342 8732 3650 8741
rect 3342 8730 3348 8732
rect 3404 8730 3428 8732
rect 3484 8730 3508 8732
rect 3564 8730 3588 8732
rect 3644 8730 3650 8732
rect 3404 8678 3406 8730
rect 3586 8678 3588 8730
rect 3342 8676 3348 8678
rect 3404 8676 3428 8678
rect 3484 8676 3508 8678
rect 3564 8676 3588 8678
rect 3644 8676 3650 8678
rect 3342 8667 3650 8676
rect 4814 8732 5122 8741
rect 4814 8730 4820 8732
rect 4876 8730 4900 8732
rect 4956 8730 4980 8732
rect 5036 8730 5060 8732
rect 5116 8730 5122 8732
rect 4876 8678 4878 8730
rect 5058 8678 5060 8730
rect 4814 8676 4820 8678
rect 4876 8676 4900 8678
rect 4956 8676 4980 8678
rect 5036 8676 5060 8678
rect 5116 8676 5122 8678
rect 4814 8667 5122 8676
rect 6286 8732 6594 8741
rect 6286 8730 6292 8732
rect 6348 8730 6372 8732
rect 6428 8730 6452 8732
rect 6508 8730 6532 8732
rect 6588 8730 6594 8732
rect 6348 8678 6350 8730
rect 6530 8678 6532 8730
rect 6286 8676 6292 8678
rect 6348 8676 6372 8678
rect 6428 8676 6452 8678
rect 6508 8676 6532 8678
rect 6588 8676 6594 8678
rect 6286 8667 6594 8676
rect 2606 8188 2914 8197
rect 2606 8186 2612 8188
rect 2668 8186 2692 8188
rect 2748 8186 2772 8188
rect 2828 8186 2852 8188
rect 2908 8186 2914 8188
rect 2668 8134 2670 8186
rect 2850 8134 2852 8186
rect 2606 8132 2612 8134
rect 2668 8132 2692 8134
rect 2748 8132 2772 8134
rect 2828 8132 2852 8134
rect 2908 8132 2914 8134
rect 2606 8123 2914 8132
rect 4078 8188 4386 8197
rect 4078 8186 4084 8188
rect 4140 8186 4164 8188
rect 4220 8186 4244 8188
rect 4300 8186 4324 8188
rect 4380 8186 4386 8188
rect 4140 8134 4142 8186
rect 4322 8134 4324 8186
rect 4078 8132 4084 8134
rect 4140 8132 4164 8134
rect 4220 8132 4244 8134
rect 4300 8132 4324 8134
rect 4380 8132 4386 8134
rect 4078 8123 4386 8132
rect 5550 8188 5858 8197
rect 5550 8186 5556 8188
rect 5612 8186 5636 8188
rect 5692 8186 5716 8188
rect 5772 8186 5796 8188
rect 5852 8186 5858 8188
rect 5612 8134 5614 8186
rect 5794 8134 5796 8186
rect 5550 8132 5556 8134
rect 5612 8132 5636 8134
rect 5692 8132 5716 8134
rect 5772 8132 5796 8134
rect 5852 8132 5858 8134
rect 5550 8123 5858 8132
rect 3342 7644 3650 7653
rect 3342 7642 3348 7644
rect 3404 7642 3428 7644
rect 3484 7642 3508 7644
rect 3564 7642 3588 7644
rect 3644 7642 3650 7644
rect 3404 7590 3406 7642
rect 3586 7590 3588 7642
rect 3342 7588 3348 7590
rect 3404 7588 3428 7590
rect 3484 7588 3508 7590
rect 3564 7588 3588 7590
rect 3644 7588 3650 7590
rect 3342 7579 3650 7588
rect 4814 7644 5122 7653
rect 4814 7642 4820 7644
rect 4876 7642 4900 7644
rect 4956 7642 4980 7644
rect 5036 7642 5060 7644
rect 5116 7642 5122 7644
rect 4876 7590 4878 7642
rect 5058 7590 5060 7642
rect 4814 7588 4820 7590
rect 4876 7588 4900 7590
rect 4956 7588 4980 7590
rect 5036 7588 5060 7590
rect 5116 7588 5122 7590
rect 4814 7579 5122 7588
rect 6286 7644 6594 7653
rect 6286 7642 6292 7644
rect 6348 7642 6372 7644
rect 6428 7642 6452 7644
rect 6508 7642 6532 7644
rect 6588 7642 6594 7644
rect 6348 7590 6350 7642
rect 6530 7590 6532 7642
rect 6286 7588 6292 7590
rect 6348 7588 6372 7590
rect 6428 7588 6452 7590
rect 6508 7588 6532 7590
rect 6588 7588 6594 7590
rect 6286 7579 6594 7588
rect 2606 7100 2914 7109
rect 2606 7098 2612 7100
rect 2668 7098 2692 7100
rect 2748 7098 2772 7100
rect 2828 7098 2852 7100
rect 2908 7098 2914 7100
rect 2668 7046 2670 7098
rect 2850 7046 2852 7098
rect 2606 7044 2612 7046
rect 2668 7044 2692 7046
rect 2748 7044 2772 7046
rect 2828 7044 2852 7046
rect 2908 7044 2914 7046
rect 2606 7035 2914 7044
rect 4078 7100 4386 7109
rect 4078 7098 4084 7100
rect 4140 7098 4164 7100
rect 4220 7098 4244 7100
rect 4300 7098 4324 7100
rect 4380 7098 4386 7100
rect 4140 7046 4142 7098
rect 4322 7046 4324 7098
rect 4078 7044 4084 7046
rect 4140 7044 4164 7046
rect 4220 7044 4244 7046
rect 4300 7044 4324 7046
rect 4380 7044 4386 7046
rect 4078 7035 4386 7044
rect 5550 7100 5858 7109
rect 5550 7098 5556 7100
rect 5612 7098 5636 7100
rect 5692 7098 5716 7100
rect 5772 7098 5796 7100
rect 5852 7098 5858 7100
rect 5612 7046 5614 7098
rect 5794 7046 5796 7098
rect 5550 7044 5556 7046
rect 5612 7044 5636 7046
rect 5692 7044 5716 7046
rect 5772 7044 5796 7046
rect 5852 7044 5858 7046
rect 5550 7035 5858 7044
rect 6932 6662 6960 9998
rect 7300 9674 7328 10202
rect 7484 10130 7512 12786
rect 7758 11996 8066 12005
rect 7758 11994 7764 11996
rect 7820 11994 7844 11996
rect 7900 11994 7924 11996
rect 7980 11994 8004 11996
rect 8060 11994 8066 11996
rect 7820 11942 7822 11994
rect 8002 11942 8004 11994
rect 7758 11940 7764 11942
rect 7820 11940 7844 11942
rect 7900 11940 7924 11942
rect 7980 11940 8004 11942
rect 8060 11940 8066 11942
rect 7758 11931 8066 11940
rect 7758 10908 8066 10917
rect 7758 10906 7764 10908
rect 7820 10906 7844 10908
rect 7900 10906 7924 10908
rect 7980 10906 8004 10908
rect 8060 10906 8066 10908
rect 7820 10854 7822 10906
rect 8002 10854 8004 10906
rect 7758 10852 7764 10854
rect 7820 10852 7844 10854
rect 7900 10852 7924 10854
rect 7980 10852 8004 10854
rect 8060 10852 8066 10854
rect 7758 10843 8066 10852
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7470 10024 7526 10033
rect 7470 9959 7526 9968
rect 7300 9646 7420 9674
rect 7022 9276 7330 9285
rect 7022 9274 7028 9276
rect 7084 9274 7108 9276
rect 7164 9274 7188 9276
rect 7244 9274 7268 9276
rect 7324 9274 7330 9276
rect 7084 9222 7086 9274
rect 7266 9222 7268 9274
rect 7022 9220 7028 9222
rect 7084 9220 7108 9222
rect 7164 9220 7188 9222
rect 7244 9220 7268 9222
rect 7324 9220 7330 9222
rect 7022 9211 7330 9220
rect 7022 8188 7330 8197
rect 7022 8186 7028 8188
rect 7084 8186 7108 8188
rect 7164 8186 7188 8188
rect 7244 8186 7268 8188
rect 7324 8186 7330 8188
rect 7084 8134 7086 8186
rect 7266 8134 7268 8186
rect 7022 8132 7028 8134
rect 7084 8132 7108 8134
rect 7164 8132 7188 8134
rect 7244 8132 7268 8134
rect 7324 8132 7330 8134
rect 7022 8123 7330 8132
rect 7022 7100 7330 7109
rect 7022 7098 7028 7100
rect 7084 7098 7108 7100
rect 7164 7098 7188 7100
rect 7244 7098 7268 7100
rect 7324 7098 7330 7100
rect 7084 7046 7086 7098
rect 7266 7046 7268 7098
rect 7022 7044 7028 7046
rect 7084 7044 7108 7046
rect 7164 7044 7188 7046
rect 7244 7044 7268 7046
rect 7324 7044 7330 7046
rect 7022 7035 7330 7044
rect 7392 6746 7420 9646
rect 7484 9450 7512 9959
rect 7576 9586 7604 10406
rect 7758 9820 8066 9829
rect 7758 9818 7764 9820
rect 7820 9818 7844 9820
rect 7900 9818 7924 9820
rect 7980 9818 8004 9820
rect 8060 9818 8066 9820
rect 7820 9766 7822 9818
rect 8002 9766 8004 9818
rect 7758 9764 7764 9766
rect 7820 9764 7844 9766
rect 7900 9764 7924 9766
rect 7980 9764 8004 9766
rect 8060 9764 8066 9766
rect 7758 9755 8066 9764
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 7758 8732 8066 8741
rect 7758 8730 7764 8732
rect 7820 8730 7844 8732
rect 7900 8730 7924 8732
rect 7980 8730 8004 8732
rect 8060 8730 8066 8732
rect 7820 8678 7822 8730
rect 8002 8678 8004 8730
rect 7758 8676 7764 8678
rect 7820 8676 7844 8678
rect 7900 8676 7924 8678
rect 7980 8676 8004 8678
rect 8060 8676 8066 8678
rect 7758 8667 8066 8676
rect 7758 7644 8066 7653
rect 7758 7642 7764 7644
rect 7820 7642 7844 7644
rect 7900 7642 7924 7644
rect 7980 7642 8004 7644
rect 8060 7642 8066 7644
rect 7820 7590 7822 7642
rect 8002 7590 8004 7642
rect 7758 7588 7764 7590
rect 7820 7588 7844 7590
rect 7900 7588 7924 7590
rect 7980 7588 8004 7590
rect 8060 7588 8066 7590
rect 7758 7579 8066 7588
rect 7392 6718 7604 6746
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 3342 6556 3650 6565
rect 3342 6554 3348 6556
rect 3404 6554 3428 6556
rect 3484 6554 3508 6556
rect 3564 6554 3588 6556
rect 3644 6554 3650 6556
rect 3404 6502 3406 6554
rect 3586 6502 3588 6554
rect 3342 6500 3348 6502
rect 3404 6500 3428 6502
rect 3484 6500 3508 6502
rect 3564 6500 3588 6502
rect 3644 6500 3650 6502
rect 3342 6491 3650 6500
rect 4814 6556 5122 6565
rect 4814 6554 4820 6556
rect 4876 6554 4900 6556
rect 4956 6554 4980 6556
rect 5036 6554 5060 6556
rect 5116 6554 5122 6556
rect 4876 6502 4878 6554
rect 5058 6502 5060 6554
rect 4814 6500 4820 6502
rect 4876 6500 4900 6502
rect 4956 6500 4980 6502
rect 5036 6500 5060 6502
rect 5116 6500 5122 6502
rect 4814 6491 5122 6500
rect 6286 6556 6594 6565
rect 6286 6554 6292 6556
rect 6348 6554 6372 6556
rect 6428 6554 6452 6556
rect 6508 6554 6532 6556
rect 6588 6554 6594 6556
rect 6348 6502 6350 6554
rect 6530 6502 6532 6554
rect 6286 6500 6292 6502
rect 6348 6500 6372 6502
rect 6428 6500 6452 6502
rect 6508 6500 6532 6502
rect 6588 6500 6594 6502
rect 6286 6491 6594 6500
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 2606 6012 2914 6021
rect 2606 6010 2612 6012
rect 2668 6010 2692 6012
rect 2748 6010 2772 6012
rect 2828 6010 2852 6012
rect 2908 6010 2914 6012
rect 2668 5958 2670 6010
rect 2850 5958 2852 6010
rect 2606 5956 2612 5958
rect 2668 5956 2692 5958
rect 2748 5956 2772 5958
rect 2828 5956 2852 5958
rect 2908 5956 2914 5958
rect 2606 5947 2914 5956
rect 4078 6012 4386 6021
rect 4078 6010 4084 6012
rect 4140 6010 4164 6012
rect 4220 6010 4244 6012
rect 4300 6010 4324 6012
rect 4380 6010 4386 6012
rect 4140 5958 4142 6010
rect 4322 5958 4324 6010
rect 4078 5956 4084 5958
rect 4140 5956 4164 5958
rect 4220 5956 4244 5958
rect 4300 5956 4324 5958
rect 4380 5956 4386 5958
rect 4078 5947 4386 5956
rect 5550 6012 5858 6021
rect 5550 6010 5556 6012
rect 5612 6010 5636 6012
rect 5692 6010 5716 6012
rect 5772 6010 5796 6012
rect 5852 6010 5858 6012
rect 5612 5958 5614 6010
rect 5794 5958 5796 6010
rect 5550 5956 5556 5958
rect 5612 5956 5636 5958
rect 5692 5956 5716 5958
rect 5772 5956 5796 5958
rect 5852 5956 5858 5958
rect 5550 5947 5858 5956
rect 6932 5914 6960 6258
rect 7022 6012 7330 6021
rect 7022 6010 7028 6012
rect 7084 6010 7108 6012
rect 7164 6010 7188 6012
rect 7244 6010 7268 6012
rect 7324 6010 7330 6012
rect 7084 5958 7086 6010
rect 7266 5958 7268 6010
rect 7022 5956 7028 5958
rect 7084 5956 7108 5958
rect 7164 5956 7188 5958
rect 7244 5956 7268 5958
rect 7324 5956 7330 5958
rect 7022 5947 7330 5956
rect 7392 5914 7420 6598
rect 7472 6112 7524 6118
rect 7470 6080 7472 6089
rect 7524 6080 7526 6089
rect 7470 6015 7526 6024
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 3342 5468 3650 5477
rect 3342 5466 3348 5468
rect 3404 5466 3428 5468
rect 3484 5466 3508 5468
rect 3564 5466 3588 5468
rect 3644 5466 3650 5468
rect 3404 5414 3406 5466
rect 3586 5414 3588 5466
rect 3342 5412 3348 5414
rect 3404 5412 3428 5414
rect 3484 5412 3508 5414
rect 3564 5412 3588 5414
rect 3644 5412 3650 5414
rect 3342 5403 3650 5412
rect 4814 5468 5122 5477
rect 4814 5466 4820 5468
rect 4876 5466 4900 5468
rect 4956 5466 4980 5468
rect 5036 5466 5060 5468
rect 5116 5466 5122 5468
rect 4876 5414 4878 5466
rect 5058 5414 5060 5466
rect 4814 5412 4820 5414
rect 4876 5412 4900 5414
rect 4956 5412 4980 5414
rect 5036 5412 5060 5414
rect 5116 5412 5122 5414
rect 4814 5403 5122 5412
rect 6286 5468 6594 5477
rect 6286 5466 6292 5468
rect 6348 5466 6372 5468
rect 6428 5466 6452 5468
rect 6508 5466 6532 5468
rect 6588 5466 6594 5468
rect 6348 5414 6350 5466
rect 6530 5414 6532 5466
rect 6286 5412 6292 5414
rect 6348 5412 6372 5414
rect 6428 5412 6452 5414
rect 6508 5412 6532 5414
rect 6588 5412 6594 5414
rect 6286 5403 6594 5412
rect 2606 4924 2914 4933
rect 2606 4922 2612 4924
rect 2668 4922 2692 4924
rect 2748 4922 2772 4924
rect 2828 4922 2852 4924
rect 2908 4922 2914 4924
rect 2668 4870 2670 4922
rect 2850 4870 2852 4922
rect 2606 4868 2612 4870
rect 2668 4868 2692 4870
rect 2748 4868 2772 4870
rect 2828 4868 2852 4870
rect 2908 4868 2914 4870
rect 2606 4859 2914 4868
rect 4078 4924 4386 4933
rect 4078 4922 4084 4924
rect 4140 4922 4164 4924
rect 4220 4922 4244 4924
rect 4300 4922 4324 4924
rect 4380 4922 4386 4924
rect 4140 4870 4142 4922
rect 4322 4870 4324 4922
rect 4078 4868 4084 4870
rect 4140 4868 4164 4870
rect 4220 4868 4244 4870
rect 4300 4868 4324 4870
rect 4380 4868 4386 4870
rect 4078 4859 4386 4868
rect 5550 4924 5858 4933
rect 5550 4922 5556 4924
rect 5612 4922 5636 4924
rect 5692 4922 5716 4924
rect 5772 4922 5796 4924
rect 5852 4922 5858 4924
rect 5612 4870 5614 4922
rect 5794 4870 5796 4922
rect 5550 4868 5556 4870
rect 5612 4868 5636 4870
rect 5692 4868 5716 4870
rect 5772 4868 5796 4870
rect 5852 4868 5858 4870
rect 5550 4859 5858 4868
rect 7022 4924 7330 4933
rect 7022 4922 7028 4924
rect 7084 4922 7108 4924
rect 7164 4922 7188 4924
rect 7244 4922 7268 4924
rect 7324 4922 7330 4924
rect 7084 4870 7086 4922
rect 7266 4870 7268 4922
rect 7022 4868 7028 4870
rect 7084 4868 7108 4870
rect 7164 4868 7188 4870
rect 7244 4868 7268 4870
rect 7324 4868 7330 4870
rect 7022 4859 7330 4868
rect 3342 4380 3650 4389
rect 3342 4378 3348 4380
rect 3404 4378 3428 4380
rect 3484 4378 3508 4380
rect 3564 4378 3588 4380
rect 3644 4378 3650 4380
rect 3404 4326 3406 4378
rect 3586 4326 3588 4378
rect 3342 4324 3348 4326
rect 3404 4324 3428 4326
rect 3484 4324 3508 4326
rect 3564 4324 3588 4326
rect 3644 4324 3650 4326
rect 3342 4315 3650 4324
rect 4814 4380 5122 4389
rect 4814 4378 4820 4380
rect 4876 4378 4900 4380
rect 4956 4378 4980 4380
rect 5036 4378 5060 4380
rect 5116 4378 5122 4380
rect 4876 4326 4878 4378
rect 5058 4326 5060 4378
rect 4814 4324 4820 4326
rect 4876 4324 4900 4326
rect 4956 4324 4980 4326
rect 5036 4324 5060 4326
rect 5116 4324 5122 4326
rect 4814 4315 5122 4324
rect 6286 4380 6594 4389
rect 6286 4378 6292 4380
rect 6348 4378 6372 4380
rect 6428 4378 6452 4380
rect 6508 4378 6532 4380
rect 6588 4378 6594 4380
rect 6348 4326 6350 4378
rect 6530 4326 6532 4378
rect 6286 4324 6292 4326
rect 6348 4324 6372 4326
rect 6428 4324 6452 4326
rect 6508 4324 6532 4326
rect 6588 4324 6594 4326
rect 6286 4315 6594 4324
rect 2606 3836 2914 3845
rect 2606 3834 2612 3836
rect 2668 3834 2692 3836
rect 2748 3834 2772 3836
rect 2828 3834 2852 3836
rect 2908 3834 2914 3836
rect 2668 3782 2670 3834
rect 2850 3782 2852 3834
rect 2606 3780 2612 3782
rect 2668 3780 2692 3782
rect 2748 3780 2772 3782
rect 2828 3780 2852 3782
rect 2908 3780 2914 3782
rect 2606 3771 2914 3780
rect 4078 3836 4386 3845
rect 4078 3834 4084 3836
rect 4140 3834 4164 3836
rect 4220 3834 4244 3836
rect 4300 3834 4324 3836
rect 4380 3834 4386 3836
rect 4140 3782 4142 3834
rect 4322 3782 4324 3834
rect 4078 3780 4084 3782
rect 4140 3780 4164 3782
rect 4220 3780 4244 3782
rect 4300 3780 4324 3782
rect 4380 3780 4386 3782
rect 4078 3771 4386 3780
rect 5550 3836 5858 3845
rect 5550 3834 5556 3836
rect 5612 3834 5636 3836
rect 5692 3834 5716 3836
rect 5772 3834 5796 3836
rect 5852 3834 5858 3836
rect 5612 3782 5614 3834
rect 5794 3782 5796 3834
rect 5550 3780 5556 3782
rect 5612 3780 5636 3782
rect 5692 3780 5716 3782
rect 5772 3780 5796 3782
rect 5852 3780 5858 3782
rect 5550 3771 5858 3780
rect 7022 3836 7330 3845
rect 7022 3834 7028 3836
rect 7084 3834 7108 3836
rect 7164 3834 7188 3836
rect 7244 3834 7268 3836
rect 7324 3834 7330 3836
rect 7084 3782 7086 3834
rect 7266 3782 7268 3834
rect 7022 3780 7028 3782
rect 7084 3780 7108 3782
rect 7164 3780 7188 3782
rect 7244 3780 7268 3782
rect 7324 3780 7330 3782
rect 7022 3771 7330 3780
rect 7392 3534 7420 5850
rect 7576 5710 7604 6718
rect 7758 6556 8066 6565
rect 7758 6554 7764 6556
rect 7820 6554 7844 6556
rect 7900 6554 7924 6556
rect 7980 6554 8004 6556
rect 8060 6554 8066 6556
rect 7820 6502 7822 6554
rect 8002 6502 8004 6554
rect 7758 6500 7764 6502
rect 7820 6500 7844 6502
rect 7900 6500 7924 6502
rect 7980 6500 8004 6502
rect 8060 6500 8066 6502
rect 7758 6491 8066 6500
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 3342 3292 3650 3301
rect 3342 3290 3348 3292
rect 3404 3290 3428 3292
rect 3484 3290 3508 3292
rect 3564 3290 3588 3292
rect 3644 3290 3650 3292
rect 3404 3238 3406 3290
rect 3586 3238 3588 3290
rect 3342 3236 3348 3238
rect 3404 3236 3428 3238
rect 3484 3236 3508 3238
rect 3564 3236 3588 3238
rect 3644 3236 3650 3238
rect 3342 3227 3650 3236
rect 4814 3292 5122 3301
rect 4814 3290 4820 3292
rect 4876 3290 4900 3292
rect 4956 3290 4980 3292
rect 5036 3290 5060 3292
rect 5116 3290 5122 3292
rect 4876 3238 4878 3290
rect 5058 3238 5060 3290
rect 4814 3236 4820 3238
rect 4876 3236 4900 3238
rect 4956 3236 4980 3238
rect 5036 3236 5060 3238
rect 5116 3236 5122 3238
rect 4814 3227 5122 3236
rect 6286 3292 6594 3301
rect 6286 3290 6292 3292
rect 6348 3290 6372 3292
rect 6428 3290 6452 3292
rect 6508 3290 6532 3292
rect 6588 3290 6594 3292
rect 6348 3238 6350 3290
rect 6530 3238 6532 3290
rect 6286 3236 6292 3238
rect 6348 3236 6372 3238
rect 6428 3236 6452 3238
rect 6508 3236 6532 3238
rect 6588 3236 6594 3238
rect 6286 3227 6594 3236
rect 6656 3058 6684 3334
rect 7392 3126 7420 3470
rect 7576 3466 7604 5646
rect 7758 5468 8066 5477
rect 7758 5466 7764 5468
rect 7820 5466 7844 5468
rect 7900 5466 7924 5468
rect 7980 5466 8004 5468
rect 8060 5466 8066 5468
rect 7820 5414 7822 5466
rect 8002 5414 8004 5466
rect 7758 5412 7764 5414
rect 7820 5412 7844 5414
rect 7900 5412 7924 5414
rect 7980 5412 8004 5414
rect 8060 5412 8066 5414
rect 7758 5403 8066 5412
rect 7758 4380 8066 4389
rect 7758 4378 7764 4380
rect 7820 4378 7844 4380
rect 7900 4378 7924 4380
rect 7980 4378 8004 4380
rect 8060 4378 8066 4380
rect 7820 4326 7822 4378
rect 8002 4326 8004 4378
rect 7758 4324 7764 4326
rect 7820 4324 7844 4326
rect 7900 4324 7924 4326
rect 7980 4324 8004 4326
rect 8060 4324 8066 4326
rect 7758 4315 8066 4324
rect 7564 3460 7616 3466
rect 7564 3402 7616 3408
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 7576 2990 7604 3402
rect 7758 3292 8066 3301
rect 7758 3290 7764 3292
rect 7820 3290 7844 3292
rect 7900 3290 7924 3292
rect 7980 3290 8004 3292
rect 8060 3290 8066 3292
rect 7820 3238 7822 3290
rect 8002 3238 8004 3290
rect 7758 3236 7764 3238
rect 7820 3236 7844 3238
rect 7900 3236 7924 3238
rect 7980 3236 8004 3238
rect 8060 3236 8066 3238
rect 7758 3227 8066 3236
rect 7564 2984 7616 2990
rect 7564 2926 7616 2932
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 2964 2848 3016 2854
rect 2964 2790 3016 2796
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 6276 2848 6328 2854
rect 6276 2790 6328 2796
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 2606 2748 2914 2757
rect 2606 2746 2612 2748
rect 2668 2746 2692 2748
rect 2748 2746 2772 2748
rect 2828 2746 2852 2748
rect 2908 2746 2914 2748
rect 2668 2694 2670 2746
rect 2850 2694 2852 2746
rect 2606 2692 2612 2694
rect 2668 2692 2692 2694
rect 2748 2692 2772 2694
rect 2828 2692 2852 2694
rect 2908 2692 2914 2694
rect 2606 2683 2914 2692
rect 2976 2446 3004 2790
rect 3896 2446 3924 2790
rect 4078 2748 4386 2757
rect 4078 2746 4084 2748
rect 4140 2746 4164 2748
rect 4220 2746 4244 2748
rect 4300 2746 4324 2748
rect 4380 2746 4386 2748
rect 4140 2694 4142 2746
rect 4322 2694 4324 2746
rect 4078 2692 4084 2694
rect 4140 2692 4164 2694
rect 4220 2692 4244 2694
rect 4300 2692 4324 2694
rect 4380 2692 4386 2694
rect 4078 2683 4386 2692
rect 5550 2748 5858 2757
rect 5550 2746 5556 2748
rect 5612 2746 5636 2748
rect 5692 2746 5716 2748
rect 5772 2746 5796 2748
rect 5852 2746 5858 2748
rect 5612 2694 5614 2746
rect 5794 2694 5796 2746
rect 5550 2692 5556 2694
rect 5612 2692 5636 2694
rect 5692 2692 5716 2694
rect 5772 2692 5796 2694
rect 5852 2692 5858 2694
rect 5550 2683 5858 2692
rect 6288 2446 6316 2790
rect 6932 2446 6960 2790
rect 7022 2748 7330 2757
rect 7022 2746 7028 2748
rect 7084 2746 7108 2748
rect 7164 2746 7188 2748
rect 7244 2746 7268 2748
rect 7324 2746 7330 2748
rect 7084 2694 7086 2746
rect 7266 2694 7268 2746
rect 7022 2692 7028 2694
rect 7084 2692 7108 2694
rect 7164 2692 7188 2694
rect 7244 2692 7268 2694
rect 7324 2692 7330 2694
rect 7022 2683 7330 2692
rect 7392 2446 7420 2858
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 1216 2372 1268 2378
rect 1216 2314 1268 2320
rect 8668 2372 8720 2378
rect 8668 2314 8720 2320
rect 1228 400 1256 2314
rect 3700 2304 3752 2310
rect 3700 2246 3752 2252
rect 6184 2304 6236 2310
rect 8208 2304 8260 2310
rect 6184 2246 6236 2252
rect 8206 2272 8208 2281
rect 8260 2272 8262 2281
rect 3342 2204 3650 2213
rect 3342 2202 3348 2204
rect 3404 2202 3428 2204
rect 3484 2202 3508 2204
rect 3564 2202 3588 2204
rect 3644 2202 3650 2204
rect 3404 2150 3406 2202
rect 3586 2150 3588 2202
rect 3342 2148 3348 2150
rect 3404 2148 3428 2150
rect 3484 2148 3508 2150
rect 3564 2148 3588 2150
rect 3644 2148 3650 2150
rect 3342 2139 3650 2148
rect 3712 400 3740 2246
rect 4814 2204 5122 2213
rect 4814 2202 4820 2204
rect 4876 2202 4900 2204
rect 4956 2202 4980 2204
rect 5036 2202 5060 2204
rect 5116 2202 5122 2204
rect 4876 2150 4878 2202
rect 5058 2150 5060 2202
rect 4814 2148 4820 2150
rect 4876 2148 4900 2150
rect 4956 2148 4980 2150
rect 5036 2148 5060 2150
rect 5116 2148 5122 2150
rect 4814 2139 5122 2148
rect 6196 400 6224 2246
rect 6286 2204 6594 2213
rect 6286 2202 6292 2204
rect 6348 2202 6372 2204
rect 6428 2202 6452 2204
rect 6508 2202 6532 2204
rect 6588 2202 6594 2204
rect 6348 2150 6350 2202
rect 6530 2150 6532 2202
rect 6286 2148 6292 2150
rect 6348 2148 6372 2150
rect 6428 2148 6452 2150
rect 6508 2148 6532 2150
rect 6588 2148 6594 2150
rect 6286 2139 6594 2148
rect 7758 2204 8066 2213
rect 8206 2207 8262 2216
rect 7758 2202 7764 2204
rect 7820 2202 7844 2204
rect 7900 2202 7924 2204
rect 7980 2202 8004 2204
rect 8060 2202 8066 2204
rect 7820 2150 7822 2202
rect 8002 2150 8004 2202
rect 7758 2148 7764 2150
rect 7820 2148 7844 2150
rect 7900 2148 7924 2150
rect 7980 2148 8004 2150
rect 8060 2148 8066 2150
rect 7758 2139 8066 2148
rect 8680 400 8708 2314
rect 1214 0 1270 400
rect 3698 0 3754 400
rect 6182 0 6238 400
rect 8666 0 8722 400
<< via2 >>
rect 2612 13626 2668 13628
rect 2692 13626 2748 13628
rect 2772 13626 2828 13628
rect 2852 13626 2908 13628
rect 2612 13574 2658 13626
rect 2658 13574 2668 13626
rect 2692 13574 2722 13626
rect 2722 13574 2734 13626
rect 2734 13574 2748 13626
rect 2772 13574 2786 13626
rect 2786 13574 2798 13626
rect 2798 13574 2828 13626
rect 2852 13574 2862 13626
rect 2862 13574 2908 13626
rect 2612 13572 2668 13574
rect 2692 13572 2748 13574
rect 2772 13572 2828 13574
rect 2852 13572 2908 13574
rect 4084 13626 4140 13628
rect 4164 13626 4220 13628
rect 4244 13626 4300 13628
rect 4324 13626 4380 13628
rect 4084 13574 4130 13626
rect 4130 13574 4140 13626
rect 4164 13574 4194 13626
rect 4194 13574 4206 13626
rect 4206 13574 4220 13626
rect 4244 13574 4258 13626
rect 4258 13574 4270 13626
rect 4270 13574 4300 13626
rect 4324 13574 4334 13626
rect 4334 13574 4380 13626
rect 4084 13572 4140 13574
rect 4164 13572 4220 13574
rect 4244 13572 4300 13574
rect 4324 13572 4380 13574
rect 5556 13626 5612 13628
rect 5636 13626 5692 13628
rect 5716 13626 5772 13628
rect 5796 13626 5852 13628
rect 5556 13574 5602 13626
rect 5602 13574 5612 13626
rect 5636 13574 5666 13626
rect 5666 13574 5678 13626
rect 5678 13574 5692 13626
rect 5716 13574 5730 13626
rect 5730 13574 5742 13626
rect 5742 13574 5772 13626
rect 5796 13574 5806 13626
rect 5806 13574 5852 13626
rect 5556 13572 5612 13574
rect 5636 13572 5692 13574
rect 5716 13572 5772 13574
rect 5796 13572 5852 13574
rect 7028 13626 7084 13628
rect 7108 13626 7164 13628
rect 7188 13626 7244 13628
rect 7268 13626 7324 13628
rect 7028 13574 7074 13626
rect 7074 13574 7084 13626
rect 7108 13574 7138 13626
rect 7138 13574 7150 13626
rect 7150 13574 7164 13626
rect 7188 13574 7202 13626
rect 7202 13574 7214 13626
rect 7214 13574 7244 13626
rect 7268 13574 7278 13626
rect 7278 13574 7324 13626
rect 7028 13572 7084 13574
rect 7108 13572 7164 13574
rect 7188 13572 7244 13574
rect 7268 13572 7324 13574
rect 8298 13640 8354 13696
rect 3348 13082 3404 13084
rect 3428 13082 3484 13084
rect 3508 13082 3564 13084
rect 3588 13082 3644 13084
rect 3348 13030 3394 13082
rect 3394 13030 3404 13082
rect 3428 13030 3458 13082
rect 3458 13030 3470 13082
rect 3470 13030 3484 13082
rect 3508 13030 3522 13082
rect 3522 13030 3534 13082
rect 3534 13030 3564 13082
rect 3588 13030 3598 13082
rect 3598 13030 3644 13082
rect 3348 13028 3404 13030
rect 3428 13028 3484 13030
rect 3508 13028 3564 13030
rect 3588 13028 3644 13030
rect 4820 13082 4876 13084
rect 4900 13082 4956 13084
rect 4980 13082 5036 13084
rect 5060 13082 5116 13084
rect 4820 13030 4866 13082
rect 4866 13030 4876 13082
rect 4900 13030 4930 13082
rect 4930 13030 4942 13082
rect 4942 13030 4956 13082
rect 4980 13030 4994 13082
rect 4994 13030 5006 13082
rect 5006 13030 5036 13082
rect 5060 13030 5070 13082
rect 5070 13030 5116 13082
rect 4820 13028 4876 13030
rect 4900 13028 4956 13030
rect 4980 13028 5036 13030
rect 5060 13028 5116 13030
rect 6292 13082 6348 13084
rect 6372 13082 6428 13084
rect 6452 13082 6508 13084
rect 6532 13082 6588 13084
rect 6292 13030 6338 13082
rect 6338 13030 6348 13082
rect 6372 13030 6402 13082
rect 6402 13030 6414 13082
rect 6414 13030 6428 13082
rect 6452 13030 6466 13082
rect 6466 13030 6478 13082
rect 6478 13030 6508 13082
rect 6532 13030 6542 13082
rect 6542 13030 6588 13082
rect 6292 13028 6348 13030
rect 6372 13028 6428 13030
rect 6452 13028 6508 13030
rect 6532 13028 6588 13030
rect 7764 13082 7820 13084
rect 7844 13082 7900 13084
rect 7924 13082 7980 13084
rect 8004 13082 8060 13084
rect 7764 13030 7810 13082
rect 7810 13030 7820 13082
rect 7844 13030 7874 13082
rect 7874 13030 7886 13082
rect 7886 13030 7900 13082
rect 7924 13030 7938 13082
rect 7938 13030 7950 13082
rect 7950 13030 7980 13082
rect 8004 13030 8014 13082
rect 8014 13030 8060 13082
rect 7764 13028 7820 13030
rect 7844 13028 7900 13030
rect 7924 13028 7980 13030
rect 8004 13028 8060 13030
rect 2612 12538 2668 12540
rect 2692 12538 2748 12540
rect 2772 12538 2828 12540
rect 2852 12538 2908 12540
rect 2612 12486 2658 12538
rect 2658 12486 2668 12538
rect 2692 12486 2722 12538
rect 2722 12486 2734 12538
rect 2734 12486 2748 12538
rect 2772 12486 2786 12538
rect 2786 12486 2798 12538
rect 2798 12486 2828 12538
rect 2852 12486 2862 12538
rect 2862 12486 2908 12538
rect 2612 12484 2668 12486
rect 2692 12484 2748 12486
rect 2772 12484 2828 12486
rect 2852 12484 2908 12486
rect 4084 12538 4140 12540
rect 4164 12538 4220 12540
rect 4244 12538 4300 12540
rect 4324 12538 4380 12540
rect 4084 12486 4130 12538
rect 4130 12486 4140 12538
rect 4164 12486 4194 12538
rect 4194 12486 4206 12538
rect 4206 12486 4220 12538
rect 4244 12486 4258 12538
rect 4258 12486 4270 12538
rect 4270 12486 4300 12538
rect 4324 12486 4334 12538
rect 4334 12486 4380 12538
rect 4084 12484 4140 12486
rect 4164 12484 4220 12486
rect 4244 12484 4300 12486
rect 4324 12484 4380 12486
rect 5556 12538 5612 12540
rect 5636 12538 5692 12540
rect 5716 12538 5772 12540
rect 5796 12538 5852 12540
rect 5556 12486 5602 12538
rect 5602 12486 5612 12538
rect 5636 12486 5666 12538
rect 5666 12486 5678 12538
rect 5678 12486 5692 12538
rect 5716 12486 5730 12538
rect 5730 12486 5742 12538
rect 5742 12486 5772 12538
rect 5796 12486 5806 12538
rect 5806 12486 5852 12538
rect 5556 12484 5612 12486
rect 5636 12484 5692 12486
rect 5716 12484 5772 12486
rect 5796 12484 5852 12486
rect 3348 11994 3404 11996
rect 3428 11994 3484 11996
rect 3508 11994 3564 11996
rect 3588 11994 3644 11996
rect 3348 11942 3394 11994
rect 3394 11942 3404 11994
rect 3428 11942 3458 11994
rect 3458 11942 3470 11994
rect 3470 11942 3484 11994
rect 3508 11942 3522 11994
rect 3522 11942 3534 11994
rect 3534 11942 3564 11994
rect 3588 11942 3598 11994
rect 3598 11942 3644 11994
rect 3348 11940 3404 11942
rect 3428 11940 3484 11942
rect 3508 11940 3564 11942
rect 3588 11940 3644 11942
rect 4820 11994 4876 11996
rect 4900 11994 4956 11996
rect 4980 11994 5036 11996
rect 5060 11994 5116 11996
rect 4820 11942 4866 11994
rect 4866 11942 4876 11994
rect 4900 11942 4930 11994
rect 4930 11942 4942 11994
rect 4942 11942 4956 11994
rect 4980 11942 4994 11994
rect 4994 11942 5006 11994
rect 5006 11942 5036 11994
rect 5060 11942 5070 11994
rect 5070 11942 5116 11994
rect 4820 11940 4876 11942
rect 4900 11940 4956 11942
rect 4980 11940 5036 11942
rect 5060 11940 5116 11942
rect 6292 11994 6348 11996
rect 6372 11994 6428 11996
rect 6452 11994 6508 11996
rect 6532 11994 6588 11996
rect 6292 11942 6338 11994
rect 6338 11942 6348 11994
rect 6372 11942 6402 11994
rect 6402 11942 6414 11994
rect 6414 11942 6428 11994
rect 6452 11942 6466 11994
rect 6466 11942 6478 11994
rect 6478 11942 6508 11994
rect 6532 11942 6542 11994
rect 6542 11942 6588 11994
rect 6292 11940 6348 11942
rect 6372 11940 6428 11942
rect 6452 11940 6508 11942
rect 6532 11940 6588 11942
rect 2612 11450 2668 11452
rect 2692 11450 2748 11452
rect 2772 11450 2828 11452
rect 2852 11450 2908 11452
rect 2612 11398 2658 11450
rect 2658 11398 2668 11450
rect 2692 11398 2722 11450
rect 2722 11398 2734 11450
rect 2734 11398 2748 11450
rect 2772 11398 2786 11450
rect 2786 11398 2798 11450
rect 2798 11398 2828 11450
rect 2852 11398 2862 11450
rect 2862 11398 2908 11450
rect 2612 11396 2668 11398
rect 2692 11396 2748 11398
rect 2772 11396 2828 11398
rect 2852 11396 2908 11398
rect 4084 11450 4140 11452
rect 4164 11450 4220 11452
rect 4244 11450 4300 11452
rect 4324 11450 4380 11452
rect 4084 11398 4130 11450
rect 4130 11398 4140 11450
rect 4164 11398 4194 11450
rect 4194 11398 4206 11450
rect 4206 11398 4220 11450
rect 4244 11398 4258 11450
rect 4258 11398 4270 11450
rect 4270 11398 4300 11450
rect 4324 11398 4334 11450
rect 4334 11398 4380 11450
rect 4084 11396 4140 11398
rect 4164 11396 4220 11398
rect 4244 11396 4300 11398
rect 4324 11396 4380 11398
rect 5556 11450 5612 11452
rect 5636 11450 5692 11452
rect 5716 11450 5772 11452
rect 5796 11450 5852 11452
rect 5556 11398 5602 11450
rect 5602 11398 5612 11450
rect 5636 11398 5666 11450
rect 5666 11398 5678 11450
rect 5678 11398 5692 11450
rect 5716 11398 5730 11450
rect 5730 11398 5742 11450
rect 5742 11398 5772 11450
rect 5796 11398 5806 11450
rect 5806 11398 5852 11450
rect 5556 11396 5612 11398
rect 5636 11396 5692 11398
rect 5716 11396 5772 11398
rect 5796 11396 5852 11398
rect 3348 10906 3404 10908
rect 3428 10906 3484 10908
rect 3508 10906 3564 10908
rect 3588 10906 3644 10908
rect 3348 10854 3394 10906
rect 3394 10854 3404 10906
rect 3428 10854 3458 10906
rect 3458 10854 3470 10906
rect 3470 10854 3484 10906
rect 3508 10854 3522 10906
rect 3522 10854 3534 10906
rect 3534 10854 3564 10906
rect 3588 10854 3598 10906
rect 3598 10854 3644 10906
rect 3348 10852 3404 10854
rect 3428 10852 3484 10854
rect 3508 10852 3564 10854
rect 3588 10852 3644 10854
rect 4820 10906 4876 10908
rect 4900 10906 4956 10908
rect 4980 10906 5036 10908
rect 5060 10906 5116 10908
rect 4820 10854 4866 10906
rect 4866 10854 4876 10906
rect 4900 10854 4930 10906
rect 4930 10854 4942 10906
rect 4942 10854 4956 10906
rect 4980 10854 4994 10906
rect 4994 10854 5006 10906
rect 5006 10854 5036 10906
rect 5060 10854 5070 10906
rect 5070 10854 5116 10906
rect 4820 10852 4876 10854
rect 4900 10852 4956 10854
rect 4980 10852 5036 10854
rect 5060 10852 5116 10854
rect 6292 10906 6348 10908
rect 6372 10906 6428 10908
rect 6452 10906 6508 10908
rect 6532 10906 6588 10908
rect 6292 10854 6338 10906
rect 6338 10854 6348 10906
rect 6372 10854 6402 10906
rect 6402 10854 6414 10906
rect 6414 10854 6428 10906
rect 6452 10854 6466 10906
rect 6466 10854 6478 10906
rect 6478 10854 6508 10906
rect 6532 10854 6542 10906
rect 6542 10854 6588 10906
rect 6292 10852 6348 10854
rect 6372 10852 6428 10854
rect 6452 10852 6508 10854
rect 6532 10852 6588 10854
rect 2612 10362 2668 10364
rect 2692 10362 2748 10364
rect 2772 10362 2828 10364
rect 2852 10362 2908 10364
rect 2612 10310 2658 10362
rect 2658 10310 2668 10362
rect 2692 10310 2722 10362
rect 2722 10310 2734 10362
rect 2734 10310 2748 10362
rect 2772 10310 2786 10362
rect 2786 10310 2798 10362
rect 2798 10310 2828 10362
rect 2852 10310 2862 10362
rect 2862 10310 2908 10362
rect 2612 10308 2668 10310
rect 2692 10308 2748 10310
rect 2772 10308 2828 10310
rect 2852 10308 2908 10310
rect 4084 10362 4140 10364
rect 4164 10362 4220 10364
rect 4244 10362 4300 10364
rect 4324 10362 4380 10364
rect 4084 10310 4130 10362
rect 4130 10310 4140 10362
rect 4164 10310 4194 10362
rect 4194 10310 4206 10362
rect 4206 10310 4220 10362
rect 4244 10310 4258 10362
rect 4258 10310 4270 10362
rect 4270 10310 4300 10362
rect 4324 10310 4334 10362
rect 4334 10310 4380 10362
rect 4084 10308 4140 10310
rect 4164 10308 4220 10310
rect 4244 10308 4300 10310
rect 4324 10308 4380 10310
rect 5556 10362 5612 10364
rect 5636 10362 5692 10364
rect 5716 10362 5772 10364
rect 5796 10362 5852 10364
rect 5556 10310 5602 10362
rect 5602 10310 5612 10362
rect 5636 10310 5666 10362
rect 5666 10310 5678 10362
rect 5678 10310 5692 10362
rect 5716 10310 5730 10362
rect 5730 10310 5742 10362
rect 5742 10310 5772 10362
rect 5796 10310 5806 10362
rect 5806 10310 5852 10362
rect 5556 10308 5612 10310
rect 5636 10308 5692 10310
rect 5716 10308 5772 10310
rect 5796 10308 5852 10310
rect 7028 12538 7084 12540
rect 7108 12538 7164 12540
rect 7188 12538 7244 12540
rect 7268 12538 7324 12540
rect 7028 12486 7074 12538
rect 7074 12486 7084 12538
rect 7108 12486 7138 12538
rect 7138 12486 7150 12538
rect 7150 12486 7164 12538
rect 7188 12486 7202 12538
rect 7202 12486 7214 12538
rect 7214 12486 7244 12538
rect 7268 12486 7278 12538
rect 7278 12486 7324 12538
rect 7028 12484 7084 12486
rect 7108 12484 7164 12486
rect 7188 12484 7244 12486
rect 7268 12484 7324 12486
rect 7028 11450 7084 11452
rect 7108 11450 7164 11452
rect 7188 11450 7244 11452
rect 7268 11450 7324 11452
rect 7028 11398 7074 11450
rect 7074 11398 7084 11450
rect 7108 11398 7138 11450
rect 7138 11398 7150 11450
rect 7150 11398 7164 11450
rect 7188 11398 7202 11450
rect 7202 11398 7214 11450
rect 7214 11398 7244 11450
rect 7268 11398 7278 11450
rect 7278 11398 7324 11450
rect 7028 11396 7084 11398
rect 7108 11396 7164 11398
rect 7188 11396 7244 11398
rect 7268 11396 7324 11398
rect 7028 10362 7084 10364
rect 7108 10362 7164 10364
rect 7188 10362 7244 10364
rect 7268 10362 7324 10364
rect 7028 10310 7074 10362
rect 7074 10310 7084 10362
rect 7108 10310 7138 10362
rect 7138 10310 7150 10362
rect 7150 10310 7164 10362
rect 7188 10310 7202 10362
rect 7202 10310 7214 10362
rect 7214 10310 7244 10362
rect 7268 10310 7278 10362
rect 7278 10310 7324 10362
rect 7028 10308 7084 10310
rect 7108 10308 7164 10310
rect 7188 10308 7244 10310
rect 7268 10308 7324 10310
rect 3348 9818 3404 9820
rect 3428 9818 3484 9820
rect 3508 9818 3564 9820
rect 3588 9818 3644 9820
rect 3348 9766 3394 9818
rect 3394 9766 3404 9818
rect 3428 9766 3458 9818
rect 3458 9766 3470 9818
rect 3470 9766 3484 9818
rect 3508 9766 3522 9818
rect 3522 9766 3534 9818
rect 3534 9766 3564 9818
rect 3588 9766 3598 9818
rect 3598 9766 3644 9818
rect 3348 9764 3404 9766
rect 3428 9764 3484 9766
rect 3508 9764 3564 9766
rect 3588 9764 3644 9766
rect 4820 9818 4876 9820
rect 4900 9818 4956 9820
rect 4980 9818 5036 9820
rect 5060 9818 5116 9820
rect 4820 9766 4866 9818
rect 4866 9766 4876 9818
rect 4900 9766 4930 9818
rect 4930 9766 4942 9818
rect 4942 9766 4956 9818
rect 4980 9766 4994 9818
rect 4994 9766 5006 9818
rect 5006 9766 5036 9818
rect 5060 9766 5070 9818
rect 5070 9766 5116 9818
rect 4820 9764 4876 9766
rect 4900 9764 4956 9766
rect 4980 9764 5036 9766
rect 5060 9764 5116 9766
rect 6292 9818 6348 9820
rect 6372 9818 6428 9820
rect 6452 9818 6508 9820
rect 6532 9818 6588 9820
rect 6292 9766 6338 9818
rect 6338 9766 6348 9818
rect 6372 9766 6402 9818
rect 6402 9766 6414 9818
rect 6414 9766 6428 9818
rect 6452 9766 6466 9818
rect 6466 9766 6478 9818
rect 6478 9766 6508 9818
rect 6532 9766 6542 9818
rect 6542 9766 6588 9818
rect 6292 9764 6348 9766
rect 6372 9764 6428 9766
rect 6452 9764 6508 9766
rect 6532 9764 6588 9766
rect 2612 9274 2668 9276
rect 2692 9274 2748 9276
rect 2772 9274 2828 9276
rect 2852 9274 2908 9276
rect 2612 9222 2658 9274
rect 2658 9222 2668 9274
rect 2692 9222 2722 9274
rect 2722 9222 2734 9274
rect 2734 9222 2748 9274
rect 2772 9222 2786 9274
rect 2786 9222 2798 9274
rect 2798 9222 2828 9274
rect 2852 9222 2862 9274
rect 2862 9222 2908 9274
rect 2612 9220 2668 9222
rect 2692 9220 2748 9222
rect 2772 9220 2828 9222
rect 2852 9220 2908 9222
rect 4084 9274 4140 9276
rect 4164 9274 4220 9276
rect 4244 9274 4300 9276
rect 4324 9274 4380 9276
rect 4084 9222 4130 9274
rect 4130 9222 4140 9274
rect 4164 9222 4194 9274
rect 4194 9222 4206 9274
rect 4206 9222 4220 9274
rect 4244 9222 4258 9274
rect 4258 9222 4270 9274
rect 4270 9222 4300 9274
rect 4324 9222 4334 9274
rect 4334 9222 4380 9274
rect 4084 9220 4140 9222
rect 4164 9220 4220 9222
rect 4244 9220 4300 9222
rect 4324 9220 4380 9222
rect 5556 9274 5612 9276
rect 5636 9274 5692 9276
rect 5716 9274 5772 9276
rect 5796 9274 5852 9276
rect 5556 9222 5602 9274
rect 5602 9222 5612 9274
rect 5636 9222 5666 9274
rect 5666 9222 5678 9274
rect 5678 9222 5692 9274
rect 5716 9222 5730 9274
rect 5730 9222 5742 9274
rect 5742 9222 5772 9274
rect 5796 9222 5806 9274
rect 5806 9222 5852 9274
rect 5556 9220 5612 9222
rect 5636 9220 5692 9222
rect 5716 9220 5772 9222
rect 5796 9220 5852 9222
rect 3348 8730 3404 8732
rect 3428 8730 3484 8732
rect 3508 8730 3564 8732
rect 3588 8730 3644 8732
rect 3348 8678 3394 8730
rect 3394 8678 3404 8730
rect 3428 8678 3458 8730
rect 3458 8678 3470 8730
rect 3470 8678 3484 8730
rect 3508 8678 3522 8730
rect 3522 8678 3534 8730
rect 3534 8678 3564 8730
rect 3588 8678 3598 8730
rect 3598 8678 3644 8730
rect 3348 8676 3404 8678
rect 3428 8676 3484 8678
rect 3508 8676 3564 8678
rect 3588 8676 3644 8678
rect 4820 8730 4876 8732
rect 4900 8730 4956 8732
rect 4980 8730 5036 8732
rect 5060 8730 5116 8732
rect 4820 8678 4866 8730
rect 4866 8678 4876 8730
rect 4900 8678 4930 8730
rect 4930 8678 4942 8730
rect 4942 8678 4956 8730
rect 4980 8678 4994 8730
rect 4994 8678 5006 8730
rect 5006 8678 5036 8730
rect 5060 8678 5070 8730
rect 5070 8678 5116 8730
rect 4820 8676 4876 8678
rect 4900 8676 4956 8678
rect 4980 8676 5036 8678
rect 5060 8676 5116 8678
rect 6292 8730 6348 8732
rect 6372 8730 6428 8732
rect 6452 8730 6508 8732
rect 6532 8730 6588 8732
rect 6292 8678 6338 8730
rect 6338 8678 6348 8730
rect 6372 8678 6402 8730
rect 6402 8678 6414 8730
rect 6414 8678 6428 8730
rect 6452 8678 6466 8730
rect 6466 8678 6478 8730
rect 6478 8678 6508 8730
rect 6532 8678 6542 8730
rect 6542 8678 6588 8730
rect 6292 8676 6348 8678
rect 6372 8676 6428 8678
rect 6452 8676 6508 8678
rect 6532 8676 6588 8678
rect 2612 8186 2668 8188
rect 2692 8186 2748 8188
rect 2772 8186 2828 8188
rect 2852 8186 2908 8188
rect 2612 8134 2658 8186
rect 2658 8134 2668 8186
rect 2692 8134 2722 8186
rect 2722 8134 2734 8186
rect 2734 8134 2748 8186
rect 2772 8134 2786 8186
rect 2786 8134 2798 8186
rect 2798 8134 2828 8186
rect 2852 8134 2862 8186
rect 2862 8134 2908 8186
rect 2612 8132 2668 8134
rect 2692 8132 2748 8134
rect 2772 8132 2828 8134
rect 2852 8132 2908 8134
rect 4084 8186 4140 8188
rect 4164 8186 4220 8188
rect 4244 8186 4300 8188
rect 4324 8186 4380 8188
rect 4084 8134 4130 8186
rect 4130 8134 4140 8186
rect 4164 8134 4194 8186
rect 4194 8134 4206 8186
rect 4206 8134 4220 8186
rect 4244 8134 4258 8186
rect 4258 8134 4270 8186
rect 4270 8134 4300 8186
rect 4324 8134 4334 8186
rect 4334 8134 4380 8186
rect 4084 8132 4140 8134
rect 4164 8132 4220 8134
rect 4244 8132 4300 8134
rect 4324 8132 4380 8134
rect 5556 8186 5612 8188
rect 5636 8186 5692 8188
rect 5716 8186 5772 8188
rect 5796 8186 5852 8188
rect 5556 8134 5602 8186
rect 5602 8134 5612 8186
rect 5636 8134 5666 8186
rect 5666 8134 5678 8186
rect 5678 8134 5692 8186
rect 5716 8134 5730 8186
rect 5730 8134 5742 8186
rect 5742 8134 5772 8186
rect 5796 8134 5806 8186
rect 5806 8134 5852 8186
rect 5556 8132 5612 8134
rect 5636 8132 5692 8134
rect 5716 8132 5772 8134
rect 5796 8132 5852 8134
rect 3348 7642 3404 7644
rect 3428 7642 3484 7644
rect 3508 7642 3564 7644
rect 3588 7642 3644 7644
rect 3348 7590 3394 7642
rect 3394 7590 3404 7642
rect 3428 7590 3458 7642
rect 3458 7590 3470 7642
rect 3470 7590 3484 7642
rect 3508 7590 3522 7642
rect 3522 7590 3534 7642
rect 3534 7590 3564 7642
rect 3588 7590 3598 7642
rect 3598 7590 3644 7642
rect 3348 7588 3404 7590
rect 3428 7588 3484 7590
rect 3508 7588 3564 7590
rect 3588 7588 3644 7590
rect 4820 7642 4876 7644
rect 4900 7642 4956 7644
rect 4980 7642 5036 7644
rect 5060 7642 5116 7644
rect 4820 7590 4866 7642
rect 4866 7590 4876 7642
rect 4900 7590 4930 7642
rect 4930 7590 4942 7642
rect 4942 7590 4956 7642
rect 4980 7590 4994 7642
rect 4994 7590 5006 7642
rect 5006 7590 5036 7642
rect 5060 7590 5070 7642
rect 5070 7590 5116 7642
rect 4820 7588 4876 7590
rect 4900 7588 4956 7590
rect 4980 7588 5036 7590
rect 5060 7588 5116 7590
rect 6292 7642 6348 7644
rect 6372 7642 6428 7644
rect 6452 7642 6508 7644
rect 6532 7642 6588 7644
rect 6292 7590 6338 7642
rect 6338 7590 6348 7642
rect 6372 7590 6402 7642
rect 6402 7590 6414 7642
rect 6414 7590 6428 7642
rect 6452 7590 6466 7642
rect 6466 7590 6478 7642
rect 6478 7590 6508 7642
rect 6532 7590 6542 7642
rect 6542 7590 6588 7642
rect 6292 7588 6348 7590
rect 6372 7588 6428 7590
rect 6452 7588 6508 7590
rect 6532 7588 6588 7590
rect 2612 7098 2668 7100
rect 2692 7098 2748 7100
rect 2772 7098 2828 7100
rect 2852 7098 2908 7100
rect 2612 7046 2658 7098
rect 2658 7046 2668 7098
rect 2692 7046 2722 7098
rect 2722 7046 2734 7098
rect 2734 7046 2748 7098
rect 2772 7046 2786 7098
rect 2786 7046 2798 7098
rect 2798 7046 2828 7098
rect 2852 7046 2862 7098
rect 2862 7046 2908 7098
rect 2612 7044 2668 7046
rect 2692 7044 2748 7046
rect 2772 7044 2828 7046
rect 2852 7044 2908 7046
rect 4084 7098 4140 7100
rect 4164 7098 4220 7100
rect 4244 7098 4300 7100
rect 4324 7098 4380 7100
rect 4084 7046 4130 7098
rect 4130 7046 4140 7098
rect 4164 7046 4194 7098
rect 4194 7046 4206 7098
rect 4206 7046 4220 7098
rect 4244 7046 4258 7098
rect 4258 7046 4270 7098
rect 4270 7046 4300 7098
rect 4324 7046 4334 7098
rect 4334 7046 4380 7098
rect 4084 7044 4140 7046
rect 4164 7044 4220 7046
rect 4244 7044 4300 7046
rect 4324 7044 4380 7046
rect 5556 7098 5612 7100
rect 5636 7098 5692 7100
rect 5716 7098 5772 7100
rect 5796 7098 5852 7100
rect 5556 7046 5602 7098
rect 5602 7046 5612 7098
rect 5636 7046 5666 7098
rect 5666 7046 5678 7098
rect 5678 7046 5692 7098
rect 5716 7046 5730 7098
rect 5730 7046 5742 7098
rect 5742 7046 5772 7098
rect 5796 7046 5806 7098
rect 5806 7046 5852 7098
rect 5556 7044 5612 7046
rect 5636 7044 5692 7046
rect 5716 7044 5772 7046
rect 5796 7044 5852 7046
rect 7764 11994 7820 11996
rect 7844 11994 7900 11996
rect 7924 11994 7980 11996
rect 8004 11994 8060 11996
rect 7764 11942 7810 11994
rect 7810 11942 7820 11994
rect 7844 11942 7874 11994
rect 7874 11942 7886 11994
rect 7886 11942 7900 11994
rect 7924 11942 7938 11994
rect 7938 11942 7950 11994
rect 7950 11942 7980 11994
rect 8004 11942 8014 11994
rect 8014 11942 8060 11994
rect 7764 11940 7820 11942
rect 7844 11940 7900 11942
rect 7924 11940 7980 11942
rect 8004 11940 8060 11942
rect 7764 10906 7820 10908
rect 7844 10906 7900 10908
rect 7924 10906 7980 10908
rect 8004 10906 8060 10908
rect 7764 10854 7810 10906
rect 7810 10854 7820 10906
rect 7844 10854 7874 10906
rect 7874 10854 7886 10906
rect 7886 10854 7900 10906
rect 7924 10854 7938 10906
rect 7938 10854 7950 10906
rect 7950 10854 7980 10906
rect 8004 10854 8014 10906
rect 8014 10854 8060 10906
rect 7764 10852 7820 10854
rect 7844 10852 7900 10854
rect 7924 10852 7980 10854
rect 8004 10852 8060 10854
rect 7470 9968 7526 10024
rect 7028 9274 7084 9276
rect 7108 9274 7164 9276
rect 7188 9274 7244 9276
rect 7268 9274 7324 9276
rect 7028 9222 7074 9274
rect 7074 9222 7084 9274
rect 7108 9222 7138 9274
rect 7138 9222 7150 9274
rect 7150 9222 7164 9274
rect 7188 9222 7202 9274
rect 7202 9222 7214 9274
rect 7214 9222 7244 9274
rect 7268 9222 7278 9274
rect 7278 9222 7324 9274
rect 7028 9220 7084 9222
rect 7108 9220 7164 9222
rect 7188 9220 7244 9222
rect 7268 9220 7324 9222
rect 7028 8186 7084 8188
rect 7108 8186 7164 8188
rect 7188 8186 7244 8188
rect 7268 8186 7324 8188
rect 7028 8134 7074 8186
rect 7074 8134 7084 8186
rect 7108 8134 7138 8186
rect 7138 8134 7150 8186
rect 7150 8134 7164 8186
rect 7188 8134 7202 8186
rect 7202 8134 7214 8186
rect 7214 8134 7244 8186
rect 7268 8134 7278 8186
rect 7278 8134 7324 8186
rect 7028 8132 7084 8134
rect 7108 8132 7164 8134
rect 7188 8132 7244 8134
rect 7268 8132 7324 8134
rect 7028 7098 7084 7100
rect 7108 7098 7164 7100
rect 7188 7098 7244 7100
rect 7268 7098 7324 7100
rect 7028 7046 7074 7098
rect 7074 7046 7084 7098
rect 7108 7046 7138 7098
rect 7138 7046 7150 7098
rect 7150 7046 7164 7098
rect 7188 7046 7202 7098
rect 7202 7046 7214 7098
rect 7214 7046 7244 7098
rect 7268 7046 7278 7098
rect 7278 7046 7324 7098
rect 7028 7044 7084 7046
rect 7108 7044 7164 7046
rect 7188 7044 7244 7046
rect 7268 7044 7324 7046
rect 7764 9818 7820 9820
rect 7844 9818 7900 9820
rect 7924 9818 7980 9820
rect 8004 9818 8060 9820
rect 7764 9766 7810 9818
rect 7810 9766 7820 9818
rect 7844 9766 7874 9818
rect 7874 9766 7886 9818
rect 7886 9766 7900 9818
rect 7924 9766 7938 9818
rect 7938 9766 7950 9818
rect 7950 9766 7980 9818
rect 8004 9766 8014 9818
rect 8014 9766 8060 9818
rect 7764 9764 7820 9766
rect 7844 9764 7900 9766
rect 7924 9764 7980 9766
rect 8004 9764 8060 9766
rect 7764 8730 7820 8732
rect 7844 8730 7900 8732
rect 7924 8730 7980 8732
rect 8004 8730 8060 8732
rect 7764 8678 7810 8730
rect 7810 8678 7820 8730
rect 7844 8678 7874 8730
rect 7874 8678 7886 8730
rect 7886 8678 7900 8730
rect 7924 8678 7938 8730
rect 7938 8678 7950 8730
rect 7950 8678 7980 8730
rect 8004 8678 8014 8730
rect 8014 8678 8060 8730
rect 7764 8676 7820 8678
rect 7844 8676 7900 8678
rect 7924 8676 7980 8678
rect 8004 8676 8060 8678
rect 7764 7642 7820 7644
rect 7844 7642 7900 7644
rect 7924 7642 7980 7644
rect 8004 7642 8060 7644
rect 7764 7590 7810 7642
rect 7810 7590 7820 7642
rect 7844 7590 7874 7642
rect 7874 7590 7886 7642
rect 7886 7590 7900 7642
rect 7924 7590 7938 7642
rect 7938 7590 7950 7642
rect 7950 7590 7980 7642
rect 8004 7590 8014 7642
rect 8014 7590 8060 7642
rect 7764 7588 7820 7590
rect 7844 7588 7900 7590
rect 7924 7588 7980 7590
rect 8004 7588 8060 7590
rect 3348 6554 3404 6556
rect 3428 6554 3484 6556
rect 3508 6554 3564 6556
rect 3588 6554 3644 6556
rect 3348 6502 3394 6554
rect 3394 6502 3404 6554
rect 3428 6502 3458 6554
rect 3458 6502 3470 6554
rect 3470 6502 3484 6554
rect 3508 6502 3522 6554
rect 3522 6502 3534 6554
rect 3534 6502 3564 6554
rect 3588 6502 3598 6554
rect 3598 6502 3644 6554
rect 3348 6500 3404 6502
rect 3428 6500 3484 6502
rect 3508 6500 3564 6502
rect 3588 6500 3644 6502
rect 4820 6554 4876 6556
rect 4900 6554 4956 6556
rect 4980 6554 5036 6556
rect 5060 6554 5116 6556
rect 4820 6502 4866 6554
rect 4866 6502 4876 6554
rect 4900 6502 4930 6554
rect 4930 6502 4942 6554
rect 4942 6502 4956 6554
rect 4980 6502 4994 6554
rect 4994 6502 5006 6554
rect 5006 6502 5036 6554
rect 5060 6502 5070 6554
rect 5070 6502 5116 6554
rect 4820 6500 4876 6502
rect 4900 6500 4956 6502
rect 4980 6500 5036 6502
rect 5060 6500 5116 6502
rect 6292 6554 6348 6556
rect 6372 6554 6428 6556
rect 6452 6554 6508 6556
rect 6532 6554 6588 6556
rect 6292 6502 6338 6554
rect 6338 6502 6348 6554
rect 6372 6502 6402 6554
rect 6402 6502 6414 6554
rect 6414 6502 6428 6554
rect 6452 6502 6466 6554
rect 6466 6502 6478 6554
rect 6478 6502 6508 6554
rect 6532 6502 6542 6554
rect 6542 6502 6588 6554
rect 6292 6500 6348 6502
rect 6372 6500 6428 6502
rect 6452 6500 6508 6502
rect 6532 6500 6588 6502
rect 2612 6010 2668 6012
rect 2692 6010 2748 6012
rect 2772 6010 2828 6012
rect 2852 6010 2908 6012
rect 2612 5958 2658 6010
rect 2658 5958 2668 6010
rect 2692 5958 2722 6010
rect 2722 5958 2734 6010
rect 2734 5958 2748 6010
rect 2772 5958 2786 6010
rect 2786 5958 2798 6010
rect 2798 5958 2828 6010
rect 2852 5958 2862 6010
rect 2862 5958 2908 6010
rect 2612 5956 2668 5958
rect 2692 5956 2748 5958
rect 2772 5956 2828 5958
rect 2852 5956 2908 5958
rect 4084 6010 4140 6012
rect 4164 6010 4220 6012
rect 4244 6010 4300 6012
rect 4324 6010 4380 6012
rect 4084 5958 4130 6010
rect 4130 5958 4140 6010
rect 4164 5958 4194 6010
rect 4194 5958 4206 6010
rect 4206 5958 4220 6010
rect 4244 5958 4258 6010
rect 4258 5958 4270 6010
rect 4270 5958 4300 6010
rect 4324 5958 4334 6010
rect 4334 5958 4380 6010
rect 4084 5956 4140 5958
rect 4164 5956 4220 5958
rect 4244 5956 4300 5958
rect 4324 5956 4380 5958
rect 5556 6010 5612 6012
rect 5636 6010 5692 6012
rect 5716 6010 5772 6012
rect 5796 6010 5852 6012
rect 5556 5958 5602 6010
rect 5602 5958 5612 6010
rect 5636 5958 5666 6010
rect 5666 5958 5678 6010
rect 5678 5958 5692 6010
rect 5716 5958 5730 6010
rect 5730 5958 5742 6010
rect 5742 5958 5772 6010
rect 5796 5958 5806 6010
rect 5806 5958 5852 6010
rect 5556 5956 5612 5958
rect 5636 5956 5692 5958
rect 5716 5956 5772 5958
rect 5796 5956 5852 5958
rect 7028 6010 7084 6012
rect 7108 6010 7164 6012
rect 7188 6010 7244 6012
rect 7268 6010 7324 6012
rect 7028 5958 7074 6010
rect 7074 5958 7084 6010
rect 7108 5958 7138 6010
rect 7138 5958 7150 6010
rect 7150 5958 7164 6010
rect 7188 5958 7202 6010
rect 7202 5958 7214 6010
rect 7214 5958 7244 6010
rect 7268 5958 7278 6010
rect 7278 5958 7324 6010
rect 7028 5956 7084 5958
rect 7108 5956 7164 5958
rect 7188 5956 7244 5958
rect 7268 5956 7324 5958
rect 7470 6060 7472 6080
rect 7472 6060 7524 6080
rect 7524 6060 7526 6080
rect 7470 6024 7526 6060
rect 3348 5466 3404 5468
rect 3428 5466 3484 5468
rect 3508 5466 3564 5468
rect 3588 5466 3644 5468
rect 3348 5414 3394 5466
rect 3394 5414 3404 5466
rect 3428 5414 3458 5466
rect 3458 5414 3470 5466
rect 3470 5414 3484 5466
rect 3508 5414 3522 5466
rect 3522 5414 3534 5466
rect 3534 5414 3564 5466
rect 3588 5414 3598 5466
rect 3598 5414 3644 5466
rect 3348 5412 3404 5414
rect 3428 5412 3484 5414
rect 3508 5412 3564 5414
rect 3588 5412 3644 5414
rect 4820 5466 4876 5468
rect 4900 5466 4956 5468
rect 4980 5466 5036 5468
rect 5060 5466 5116 5468
rect 4820 5414 4866 5466
rect 4866 5414 4876 5466
rect 4900 5414 4930 5466
rect 4930 5414 4942 5466
rect 4942 5414 4956 5466
rect 4980 5414 4994 5466
rect 4994 5414 5006 5466
rect 5006 5414 5036 5466
rect 5060 5414 5070 5466
rect 5070 5414 5116 5466
rect 4820 5412 4876 5414
rect 4900 5412 4956 5414
rect 4980 5412 5036 5414
rect 5060 5412 5116 5414
rect 6292 5466 6348 5468
rect 6372 5466 6428 5468
rect 6452 5466 6508 5468
rect 6532 5466 6588 5468
rect 6292 5414 6338 5466
rect 6338 5414 6348 5466
rect 6372 5414 6402 5466
rect 6402 5414 6414 5466
rect 6414 5414 6428 5466
rect 6452 5414 6466 5466
rect 6466 5414 6478 5466
rect 6478 5414 6508 5466
rect 6532 5414 6542 5466
rect 6542 5414 6588 5466
rect 6292 5412 6348 5414
rect 6372 5412 6428 5414
rect 6452 5412 6508 5414
rect 6532 5412 6588 5414
rect 2612 4922 2668 4924
rect 2692 4922 2748 4924
rect 2772 4922 2828 4924
rect 2852 4922 2908 4924
rect 2612 4870 2658 4922
rect 2658 4870 2668 4922
rect 2692 4870 2722 4922
rect 2722 4870 2734 4922
rect 2734 4870 2748 4922
rect 2772 4870 2786 4922
rect 2786 4870 2798 4922
rect 2798 4870 2828 4922
rect 2852 4870 2862 4922
rect 2862 4870 2908 4922
rect 2612 4868 2668 4870
rect 2692 4868 2748 4870
rect 2772 4868 2828 4870
rect 2852 4868 2908 4870
rect 4084 4922 4140 4924
rect 4164 4922 4220 4924
rect 4244 4922 4300 4924
rect 4324 4922 4380 4924
rect 4084 4870 4130 4922
rect 4130 4870 4140 4922
rect 4164 4870 4194 4922
rect 4194 4870 4206 4922
rect 4206 4870 4220 4922
rect 4244 4870 4258 4922
rect 4258 4870 4270 4922
rect 4270 4870 4300 4922
rect 4324 4870 4334 4922
rect 4334 4870 4380 4922
rect 4084 4868 4140 4870
rect 4164 4868 4220 4870
rect 4244 4868 4300 4870
rect 4324 4868 4380 4870
rect 5556 4922 5612 4924
rect 5636 4922 5692 4924
rect 5716 4922 5772 4924
rect 5796 4922 5852 4924
rect 5556 4870 5602 4922
rect 5602 4870 5612 4922
rect 5636 4870 5666 4922
rect 5666 4870 5678 4922
rect 5678 4870 5692 4922
rect 5716 4870 5730 4922
rect 5730 4870 5742 4922
rect 5742 4870 5772 4922
rect 5796 4870 5806 4922
rect 5806 4870 5852 4922
rect 5556 4868 5612 4870
rect 5636 4868 5692 4870
rect 5716 4868 5772 4870
rect 5796 4868 5852 4870
rect 7028 4922 7084 4924
rect 7108 4922 7164 4924
rect 7188 4922 7244 4924
rect 7268 4922 7324 4924
rect 7028 4870 7074 4922
rect 7074 4870 7084 4922
rect 7108 4870 7138 4922
rect 7138 4870 7150 4922
rect 7150 4870 7164 4922
rect 7188 4870 7202 4922
rect 7202 4870 7214 4922
rect 7214 4870 7244 4922
rect 7268 4870 7278 4922
rect 7278 4870 7324 4922
rect 7028 4868 7084 4870
rect 7108 4868 7164 4870
rect 7188 4868 7244 4870
rect 7268 4868 7324 4870
rect 3348 4378 3404 4380
rect 3428 4378 3484 4380
rect 3508 4378 3564 4380
rect 3588 4378 3644 4380
rect 3348 4326 3394 4378
rect 3394 4326 3404 4378
rect 3428 4326 3458 4378
rect 3458 4326 3470 4378
rect 3470 4326 3484 4378
rect 3508 4326 3522 4378
rect 3522 4326 3534 4378
rect 3534 4326 3564 4378
rect 3588 4326 3598 4378
rect 3598 4326 3644 4378
rect 3348 4324 3404 4326
rect 3428 4324 3484 4326
rect 3508 4324 3564 4326
rect 3588 4324 3644 4326
rect 4820 4378 4876 4380
rect 4900 4378 4956 4380
rect 4980 4378 5036 4380
rect 5060 4378 5116 4380
rect 4820 4326 4866 4378
rect 4866 4326 4876 4378
rect 4900 4326 4930 4378
rect 4930 4326 4942 4378
rect 4942 4326 4956 4378
rect 4980 4326 4994 4378
rect 4994 4326 5006 4378
rect 5006 4326 5036 4378
rect 5060 4326 5070 4378
rect 5070 4326 5116 4378
rect 4820 4324 4876 4326
rect 4900 4324 4956 4326
rect 4980 4324 5036 4326
rect 5060 4324 5116 4326
rect 6292 4378 6348 4380
rect 6372 4378 6428 4380
rect 6452 4378 6508 4380
rect 6532 4378 6588 4380
rect 6292 4326 6338 4378
rect 6338 4326 6348 4378
rect 6372 4326 6402 4378
rect 6402 4326 6414 4378
rect 6414 4326 6428 4378
rect 6452 4326 6466 4378
rect 6466 4326 6478 4378
rect 6478 4326 6508 4378
rect 6532 4326 6542 4378
rect 6542 4326 6588 4378
rect 6292 4324 6348 4326
rect 6372 4324 6428 4326
rect 6452 4324 6508 4326
rect 6532 4324 6588 4326
rect 2612 3834 2668 3836
rect 2692 3834 2748 3836
rect 2772 3834 2828 3836
rect 2852 3834 2908 3836
rect 2612 3782 2658 3834
rect 2658 3782 2668 3834
rect 2692 3782 2722 3834
rect 2722 3782 2734 3834
rect 2734 3782 2748 3834
rect 2772 3782 2786 3834
rect 2786 3782 2798 3834
rect 2798 3782 2828 3834
rect 2852 3782 2862 3834
rect 2862 3782 2908 3834
rect 2612 3780 2668 3782
rect 2692 3780 2748 3782
rect 2772 3780 2828 3782
rect 2852 3780 2908 3782
rect 4084 3834 4140 3836
rect 4164 3834 4220 3836
rect 4244 3834 4300 3836
rect 4324 3834 4380 3836
rect 4084 3782 4130 3834
rect 4130 3782 4140 3834
rect 4164 3782 4194 3834
rect 4194 3782 4206 3834
rect 4206 3782 4220 3834
rect 4244 3782 4258 3834
rect 4258 3782 4270 3834
rect 4270 3782 4300 3834
rect 4324 3782 4334 3834
rect 4334 3782 4380 3834
rect 4084 3780 4140 3782
rect 4164 3780 4220 3782
rect 4244 3780 4300 3782
rect 4324 3780 4380 3782
rect 5556 3834 5612 3836
rect 5636 3834 5692 3836
rect 5716 3834 5772 3836
rect 5796 3834 5852 3836
rect 5556 3782 5602 3834
rect 5602 3782 5612 3834
rect 5636 3782 5666 3834
rect 5666 3782 5678 3834
rect 5678 3782 5692 3834
rect 5716 3782 5730 3834
rect 5730 3782 5742 3834
rect 5742 3782 5772 3834
rect 5796 3782 5806 3834
rect 5806 3782 5852 3834
rect 5556 3780 5612 3782
rect 5636 3780 5692 3782
rect 5716 3780 5772 3782
rect 5796 3780 5852 3782
rect 7028 3834 7084 3836
rect 7108 3834 7164 3836
rect 7188 3834 7244 3836
rect 7268 3834 7324 3836
rect 7028 3782 7074 3834
rect 7074 3782 7084 3834
rect 7108 3782 7138 3834
rect 7138 3782 7150 3834
rect 7150 3782 7164 3834
rect 7188 3782 7202 3834
rect 7202 3782 7214 3834
rect 7214 3782 7244 3834
rect 7268 3782 7278 3834
rect 7278 3782 7324 3834
rect 7028 3780 7084 3782
rect 7108 3780 7164 3782
rect 7188 3780 7244 3782
rect 7268 3780 7324 3782
rect 7764 6554 7820 6556
rect 7844 6554 7900 6556
rect 7924 6554 7980 6556
rect 8004 6554 8060 6556
rect 7764 6502 7810 6554
rect 7810 6502 7820 6554
rect 7844 6502 7874 6554
rect 7874 6502 7886 6554
rect 7886 6502 7900 6554
rect 7924 6502 7938 6554
rect 7938 6502 7950 6554
rect 7950 6502 7980 6554
rect 8004 6502 8014 6554
rect 8014 6502 8060 6554
rect 7764 6500 7820 6502
rect 7844 6500 7900 6502
rect 7924 6500 7980 6502
rect 8004 6500 8060 6502
rect 3348 3290 3404 3292
rect 3428 3290 3484 3292
rect 3508 3290 3564 3292
rect 3588 3290 3644 3292
rect 3348 3238 3394 3290
rect 3394 3238 3404 3290
rect 3428 3238 3458 3290
rect 3458 3238 3470 3290
rect 3470 3238 3484 3290
rect 3508 3238 3522 3290
rect 3522 3238 3534 3290
rect 3534 3238 3564 3290
rect 3588 3238 3598 3290
rect 3598 3238 3644 3290
rect 3348 3236 3404 3238
rect 3428 3236 3484 3238
rect 3508 3236 3564 3238
rect 3588 3236 3644 3238
rect 4820 3290 4876 3292
rect 4900 3290 4956 3292
rect 4980 3290 5036 3292
rect 5060 3290 5116 3292
rect 4820 3238 4866 3290
rect 4866 3238 4876 3290
rect 4900 3238 4930 3290
rect 4930 3238 4942 3290
rect 4942 3238 4956 3290
rect 4980 3238 4994 3290
rect 4994 3238 5006 3290
rect 5006 3238 5036 3290
rect 5060 3238 5070 3290
rect 5070 3238 5116 3290
rect 4820 3236 4876 3238
rect 4900 3236 4956 3238
rect 4980 3236 5036 3238
rect 5060 3236 5116 3238
rect 6292 3290 6348 3292
rect 6372 3290 6428 3292
rect 6452 3290 6508 3292
rect 6532 3290 6588 3292
rect 6292 3238 6338 3290
rect 6338 3238 6348 3290
rect 6372 3238 6402 3290
rect 6402 3238 6414 3290
rect 6414 3238 6428 3290
rect 6452 3238 6466 3290
rect 6466 3238 6478 3290
rect 6478 3238 6508 3290
rect 6532 3238 6542 3290
rect 6542 3238 6588 3290
rect 6292 3236 6348 3238
rect 6372 3236 6428 3238
rect 6452 3236 6508 3238
rect 6532 3236 6588 3238
rect 7764 5466 7820 5468
rect 7844 5466 7900 5468
rect 7924 5466 7980 5468
rect 8004 5466 8060 5468
rect 7764 5414 7810 5466
rect 7810 5414 7820 5466
rect 7844 5414 7874 5466
rect 7874 5414 7886 5466
rect 7886 5414 7900 5466
rect 7924 5414 7938 5466
rect 7938 5414 7950 5466
rect 7950 5414 7980 5466
rect 8004 5414 8014 5466
rect 8014 5414 8060 5466
rect 7764 5412 7820 5414
rect 7844 5412 7900 5414
rect 7924 5412 7980 5414
rect 8004 5412 8060 5414
rect 7764 4378 7820 4380
rect 7844 4378 7900 4380
rect 7924 4378 7980 4380
rect 8004 4378 8060 4380
rect 7764 4326 7810 4378
rect 7810 4326 7820 4378
rect 7844 4326 7874 4378
rect 7874 4326 7886 4378
rect 7886 4326 7900 4378
rect 7924 4326 7938 4378
rect 7938 4326 7950 4378
rect 7950 4326 7980 4378
rect 8004 4326 8014 4378
rect 8014 4326 8060 4378
rect 7764 4324 7820 4326
rect 7844 4324 7900 4326
rect 7924 4324 7980 4326
rect 8004 4324 8060 4326
rect 7764 3290 7820 3292
rect 7844 3290 7900 3292
rect 7924 3290 7980 3292
rect 8004 3290 8060 3292
rect 7764 3238 7810 3290
rect 7810 3238 7820 3290
rect 7844 3238 7874 3290
rect 7874 3238 7886 3290
rect 7886 3238 7900 3290
rect 7924 3238 7938 3290
rect 7938 3238 7950 3290
rect 7950 3238 7980 3290
rect 8004 3238 8014 3290
rect 8014 3238 8060 3290
rect 7764 3236 7820 3238
rect 7844 3236 7900 3238
rect 7924 3236 7980 3238
rect 8004 3236 8060 3238
rect 2612 2746 2668 2748
rect 2692 2746 2748 2748
rect 2772 2746 2828 2748
rect 2852 2746 2908 2748
rect 2612 2694 2658 2746
rect 2658 2694 2668 2746
rect 2692 2694 2722 2746
rect 2722 2694 2734 2746
rect 2734 2694 2748 2746
rect 2772 2694 2786 2746
rect 2786 2694 2798 2746
rect 2798 2694 2828 2746
rect 2852 2694 2862 2746
rect 2862 2694 2908 2746
rect 2612 2692 2668 2694
rect 2692 2692 2748 2694
rect 2772 2692 2828 2694
rect 2852 2692 2908 2694
rect 4084 2746 4140 2748
rect 4164 2746 4220 2748
rect 4244 2746 4300 2748
rect 4324 2746 4380 2748
rect 4084 2694 4130 2746
rect 4130 2694 4140 2746
rect 4164 2694 4194 2746
rect 4194 2694 4206 2746
rect 4206 2694 4220 2746
rect 4244 2694 4258 2746
rect 4258 2694 4270 2746
rect 4270 2694 4300 2746
rect 4324 2694 4334 2746
rect 4334 2694 4380 2746
rect 4084 2692 4140 2694
rect 4164 2692 4220 2694
rect 4244 2692 4300 2694
rect 4324 2692 4380 2694
rect 5556 2746 5612 2748
rect 5636 2746 5692 2748
rect 5716 2746 5772 2748
rect 5796 2746 5852 2748
rect 5556 2694 5602 2746
rect 5602 2694 5612 2746
rect 5636 2694 5666 2746
rect 5666 2694 5678 2746
rect 5678 2694 5692 2746
rect 5716 2694 5730 2746
rect 5730 2694 5742 2746
rect 5742 2694 5772 2746
rect 5796 2694 5806 2746
rect 5806 2694 5852 2746
rect 5556 2692 5612 2694
rect 5636 2692 5692 2694
rect 5716 2692 5772 2694
rect 5796 2692 5852 2694
rect 7028 2746 7084 2748
rect 7108 2746 7164 2748
rect 7188 2746 7244 2748
rect 7268 2746 7324 2748
rect 7028 2694 7074 2746
rect 7074 2694 7084 2746
rect 7108 2694 7138 2746
rect 7138 2694 7150 2746
rect 7150 2694 7164 2746
rect 7188 2694 7202 2746
rect 7202 2694 7214 2746
rect 7214 2694 7244 2746
rect 7268 2694 7278 2746
rect 7278 2694 7324 2746
rect 7028 2692 7084 2694
rect 7108 2692 7164 2694
rect 7188 2692 7244 2694
rect 7268 2692 7324 2694
rect 8206 2252 8208 2272
rect 8208 2252 8260 2272
rect 8260 2252 8262 2272
rect 3348 2202 3404 2204
rect 3428 2202 3484 2204
rect 3508 2202 3564 2204
rect 3588 2202 3644 2204
rect 3348 2150 3394 2202
rect 3394 2150 3404 2202
rect 3428 2150 3458 2202
rect 3458 2150 3470 2202
rect 3470 2150 3484 2202
rect 3508 2150 3522 2202
rect 3522 2150 3534 2202
rect 3534 2150 3564 2202
rect 3588 2150 3598 2202
rect 3598 2150 3644 2202
rect 3348 2148 3404 2150
rect 3428 2148 3484 2150
rect 3508 2148 3564 2150
rect 3588 2148 3644 2150
rect 4820 2202 4876 2204
rect 4900 2202 4956 2204
rect 4980 2202 5036 2204
rect 5060 2202 5116 2204
rect 4820 2150 4866 2202
rect 4866 2150 4876 2202
rect 4900 2150 4930 2202
rect 4930 2150 4942 2202
rect 4942 2150 4956 2202
rect 4980 2150 4994 2202
rect 4994 2150 5006 2202
rect 5006 2150 5036 2202
rect 5060 2150 5070 2202
rect 5070 2150 5116 2202
rect 4820 2148 4876 2150
rect 4900 2148 4956 2150
rect 4980 2148 5036 2150
rect 5060 2148 5116 2150
rect 8206 2216 8262 2252
rect 6292 2202 6348 2204
rect 6372 2202 6428 2204
rect 6452 2202 6508 2204
rect 6532 2202 6588 2204
rect 6292 2150 6338 2202
rect 6338 2150 6348 2202
rect 6372 2150 6402 2202
rect 6402 2150 6414 2202
rect 6414 2150 6428 2202
rect 6452 2150 6466 2202
rect 6466 2150 6478 2202
rect 6478 2150 6508 2202
rect 6532 2150 6542 2202
rect 6542 2150 6588 2202
rect 6292 2148 6348 2150
rect 6372 2148 6428 2150
rect 6452 2148 6508 2150
rect 6532 2148 6588 2150
rect 7764 2202 7820 2204
rect 7844 2202 7900 2204
rect 7924 2202 7980 2204
rect 8004 2202 8060 2204
rect 7764 2150 7810 2202
rect 7810 2150 7820 2202
rect 7844 2150 7874 2202
rect 7874 2150 7886 2202
rect 7886 2150 7900 2202
rect 7924 2150 7938 2202
rect 7938 2150 7950 2202
rect 7950 2150 7980 2202
rect 8004 2150 8014 2202
rect 8014 2150 8060 2202
rect 7764 2148 7820 2150
rect 7844 2148 7900 2150
rect 7924 2148 7980 2150
rect 8004 2148 8060 2150
<< metal3 >>
rect 8293 13698 8359 13701
rect 9600 13698 10000 13728
rect 8293 13696 10000 13698
rect 8293 13640 8298 13696
rect 8354 13640 10000 13696
rect 8293 13638 10000 13640
rect 8293 13635 8359 13638
rect 2602 13632 2918 13633
rect 2602 13568 2608 13632
rect 2672 13568 2688 13632
rect 2752 13568 2768 13632
rect 2832 13568 2848 13632
rect 2912 13568 2918 13632
rect 2602 13567 2918 13568
rect 4074 13632 4390 13633
rect 4074 13568 4080 13632
rect 4144 13568 4160 13632
rect 4224 13568 4240 13632
rect 4304 13568 4320 13632
rect 4384 13568 4390 13632
rect 4074 13567 4390 13568
rect 5546 13632 5862 13633
rect 5546 13568 5552 13632
rect 5616 13568 5632 13632
rect 5696 13568 5712 13632
rect 5776 13568 5792 13632
rect 5856 13568 5862 13632
rect 5546 13567 5862 13568
rect 7018 13632 7334 13633
rect 7018 13568 7024 13632
rect 7088 13568 7104 13632
rect 7168 13568 7184 13632
rect 7248 13568 7264 13632
rect 7328 13568 7334 13632
rect 9600 13608 10000 13638
rect 7018 13567 7334 13568
rect 3338 13088 3654 13089
rect 3338 13024 3344 13088
rect 3408 13024 3424 13088
rect 3488 13024 3504 13088
rect 3568 13024 3584 13088
rect 3648 13024 3654 13088
rect 3338 13023 3654 13024
rect 4810 13088 5126 13089
rect 4810 13024 4816 13088
rect 4880 13024 4896 13088
rect 4960 13024 4976 13088
rect 5040 13024 5056 13088
rect 5120 13024 5126 13088
rect 4810 13023 5126 13024
rect 6282 13088 6598 13089
rect 6282 13024 6288 13088
rect 6352 13024 6368 13088
rect 6432 13024 6448 13088
rect 6512 13024 6528 13088
rect 6592 13024 6598 13088
rect 6282 13023 6598 13024
rect 7754 13088 8070 13089
rect 7754 13024 7760 13088
rect 7824 13024 7840 13088
rect 7904 13024 7920 13088
rect 7984 13024 8000 13088
rect 8064 13024 8070 13088
rect 7754 13023 8070 13024
rect 2602 12544 2918 12545
rect 2602 12480 2608 12544
rect 2672 12480 2688 12544
rect 2752 12480 2768 12544
rect 2832 12480 2848 12544
rect 2912 12480 2918 12544
rect 2602 12479 2918 12480
rect 4074 12544 4390 12545
rect 4074 12480 4080 12544
rect 4144 12480 4160 12544
rect 4224 12480 4240 12544
rect 4304 12480 4320 12544
rect 4384 12480 4390 12544
rect 4074 12479 4390 12480
rect 5546 12544 5862 12545
rect 5546 12480 5552 12544
rect 5616 12480 5632 12544
rect 5696 12480 5712 12544
rect 5776 12480 5792 12544
rect 5856 12480 5862 12544
rect 5546 12479 5862 12480
rect 7018 12544 7334 12545
rect 7018 12480 7024 12544
rect 7088 12480 7104 12544
rect 7168 12480 7184 12544
rect 7248 12480 7264 12544
rect 7328 12480 7334 12544
rect 7018 12479 7334 12480
rect 3338 12000 3654 12001
rect 3338 11936 3344 12000
rect 3408 11936 3424 12000
rect 3488 11936 3504 12000
rect 3568 11936 3584 12000
rect 3648 11936 3654 12000
rect 3338 11935 3654 11936
rect 4810 12000 5126 12001
rect 4810 11936 4816 12000
rect 4880 11936 4896 12000
rect 4960 11936 4976 12000
rect 5040 11936 5056 12000
rect 5120 11936 5126 12000
rect 4810 11935 5126 11936
rect 6282 12000 6598 12001
rect 6282 11936 6288 12000
rect 6352 11936 6368 12000
rect 6432 11936 6448 12000
rect 6512 11936 6528 12000
rect 6592 11936 6598 12000
rect 6282 11935 6598 11936
rect 7754 12000 8070 12001
rect 7754 11936 7760 12000
rect 7824 11936 7840 12000
rect 7904 11936 7920 12000
rect 7984 11936 8000 12000
rect 8064 11936 8070 12000
rect 7754 11935 8070 11936
rect 2602 11456 2918 11457
rect 2602 11392 2608 11456
rect 2672 11392 2688 11456
rect 2752 11392 2768 11456
rect 2832 11392 2848 11456
rect 2912 11392 2918 11456
rect 2602 11391 2918 11392
rect 4074 11456 4390 11457
rect 4074 11392 4080 11456
rect 4144 11392 4160 11456
rect 4224 11392 4240 11456
rect 4304 11392 4320 11456
rect 4384 11392 4390 11456
rect 4074 11391 4390 11392
rect 5546 11456 5862 11457
rect 5546 11392 5552 11456
rect 5616 11392 5632 11456
rect 5696 11392 5712 11456
rect 5776 11392 5792 11456
rect 5856 11392 5862 11456
rect 5546 11391 5862 11392
rect 7018 11456 7334 11457
rect 7018 11392 7024 11456
rect 7088 11392 7104 11456
rect 7168 11392 7184 11456
rect 7248 11392 7264 11456
rect 7328 11392 7334 11456
rect 7018 11391 7334 11392
rect 3338 10912 3654 10913
rect 3338 10848 3344 10912
rect 3408 10848 3424 10912
rect 3488 10848 3504 10912
rect 3568 10848 3584 10912
rect 3648 10848 3654 10912
rect 3338 10847 3654 10848
rect 4810 10912 5126 10913
rect 4810 10848 4816 10912
rect 4880 10848 4896 10912
rect 4960 10848 4976 10912
rect 5040 10848 5056 10912
rect 5120 10848 5126 10912
rect 4810 10847 5126 10848
rect 6282 10912 6598 10913
rect 6282 10848 6288 10912
rect 6352 10848 6368 10912
rect 6432 10848 6448 10912
rect 6512 10848 6528 10912
rect 6592 10848 6598 10912
rect 6282 10847 6598 10848
rect 7754 10912 8070 10913
rect 7754 10848 7760 10912
rect 7824 10848 7840 10912
rect 7904 10848 7920 10912
rect 7984 10848 8000 10912
rect 8064 10848 8070 10912
rect 7754 10847 8070 10848
rect 2602 10368 2918 10369
rect 2602 10304 2608 10368
rect 2672 10304 2688 10368
rect 2752 10304 2768 10368
rect 2832 10304 2848 10368
rect 2912 10304 2918 10368
rect 2602 10303 2918 10304
rect 4074 10368 4390 10369
rect 4074 10304 4080 10368
rect 4144 10304 4160 10368
rect 4224 10304 4240 10368
rect 4304 10304 4320 10368
rect 4384 10304 4390 10368
rect 4074 10303 4390 10304
rect 5546 10368 5862 10369
rect 5546 10304 5552 10368
rect 5616 10304 5632 10368
rect 5696 10304 5712 10368
rect 5776 10304 5792 10368
rect 5856 10304 5862 10368
rect 5546 10303 5862 10304
rect 7018 10368 7334 10369
rect 7018 10304 7024 10368
rect 7088 10304 7104 10368
rect 7168 10304 7184 10368
rect 7248 10304 7264 10368
rect 7328 10304 7334 10368
rect 7018 10303 7334 10304
rect 7465 10026 7531 10029
rect 7465 10024 8218 10026
rect 7465 9968 7470 10024
rect 7526 9968 8218 10024
rect 7465 9966 8218 9968
rect 7465 9963 7531 9966
rect 8158 9890 8218 9966
rect 9600 9890 10000 9920
rect 8158 9830 10000 9890
rect 3338 9824 3654 9825
rect 3338 9760 3344 9824
rect 3408 9760 3424 9824
rect 3488 9760 3504 9824
rect 3568 9760 3584 9824
rect 3648 9760 3654 9824
rect 3338 9759 3654 9760
rect 4810 9824 5126 9825
rect 4810 9760 4816 9824
rect 4880 9760 4896 9824
rect 4960 9760 4976 9824
rect 5040 9760 5056 9824
rect 5120 9760 5126 9824
rect 4810 9759 5126 9760
rect 6282 9824 6598 9825
rect 6282 9760 6288 9824
rect 6352 9760 6368 9824
rect 6432 9760 6448 9824
rect 6512 9760 6528 9824
rect 6592 9760 6598 9824
rect 6282 9759 6598 9760
rect 7754 9824 8070 9825
rect 7754 9760 7760 9824
rect 7824 9760 7840 9824
rect 7904 9760 7920 9824
rect 7984 9760 8000 9824
rect 8064 9760 8070 9824
rect 9600 9800 10000 9830
rect 7754 9759 8070 9760
rect 2602 9280 2918 9281
rect 2602 9216 2608 9280
rect 2672 9216 2688 9280
rect 2752 9216 2768 9280
rect 2832 9216 2848 9280
rect 2912 9216 2918 9280
rect 2602 9215 2918 9216
rect 4074 9280 4390 9281
rect 4074 9216 4080 9280
rect 4144 9216 4160 9280
rect 4224 9216 4240 9280
rect 4304 9216 4320 9280
rect 4384 9216 4390 9280
rect 4074 9215 4390 9216
rect 5546 9280 5862 9281
rect 5546 9216 5552 9280
rect 5616 9216 5632 9280
rect 5696 9216 5712 9280
rect 5776 9216 5792 9280
rect 5856 9216 5862 9280
rect 5546 9215 5862 9216
rect 7018 9280 7334 9281
rect 7018 9216 7024 9280
rect 7088 9216 7104 9280
rect 7168 9216 7184 9280
rect 7248 9216 7264 9280
rect 7328 9216 7334 9280
rect 7018 9215 7334 9216
rect 3338 8736 3654 8737
rect 3338 8672 3344 8736
rect 3408 8672 3424 8736
rect 3488 8672 3504 8736
rect 3568 8672 3584 8736
rect 3648 8672 3654 8736
rect 3338 8671 3654 8672
rect 4810 8736 5126 8737
rect 4810 8672 4816 8736
rect 4880 8672 4896 8736
rect 4960 8672 4976 8736
rect 5040 8672 5056 8736
rect 5120 8672 5126 8736
rect 4810 8671 5126 8672
rect 6282 8736 6598 8737
rect 6282 8672 6288 8736
rect 6352 8672 6368 8736
rect 6432 8672 6448 8736
rect 6512 8672 6528 8736
rect 6592 8672 6598 8736
rect 6282 8671 6598 8672
rect 7754 8736 8070 8737
rect 7754 8672 7760 8736
rect 7824 8672 7840 8736
rect 7904 8672 7920 8736
rect 7984 8672 8000 8736
rect 8064 8672 8070 8736
rect 7754 8671 8070 8672
rect 2602 8192 2918 8193
rect 2602 8128 2608 8192
rect 2672 8128 2688 8192
rect 2752 8128 2768 8192
rect 2832 8128 2848 8192
rect 2912 8128 2918 8192
rect 2602 8127 2918 8128
rect 4074 8192 4390 8193
rect 4074 8128 4080 8192
rect 4144 8128 4160 8192
rect 4224 8128 4240 8192
rect 4304 8128 4320 8192
rect 4384 8128 4390 8192
rect 4074 8127 4390 8128
rect 5546 8192 5862 8193
rect 5546 8128 5552 8192
rect 5616 8128 5632 8192
rect 5696 8128 5712 8192
rect 5776 8128 5792 8192
rect 5856 8128 5862 8192
rect 5546 8127 5862 8128
rect 7018 8192 7334 8193
rect 7018 8128 7024 8192
rect 7088 8128 7104 8192
rect 7168 8128 7184 8192
rect 7248 8128 7264 8192
rect 7328 8128 7334 8192
rect 7018 8127 7334 8128
rect 3338 7648 3654 7649
rect 3338 7584 3344 7648
rect 3408 7584 3424 7648
rect 3488 7584 3504 7648
rect 3568 7584 3584 7648
rect 3648 7584 3654 7648
rect 3338 7583 3654 7584
rect 4810 7648 5126 7649
rect 4810 7584 4816 7648
rect 4880 7584 4896 7648
rect 4960 7584 4976 7648
rect 5040 7584 5056 7648
rect 5120 7584 5126 7648
rect 4810 7583 5126 7584
rect 6282 7648 6598 7649
rect 6282 7584 6288 7648
rect 6352 7584 6368 7648
rect 6432 7584 6448 7648
rect 6512 7584 6528 7648
rect 6592 7584 6598 7648
rect 6282 7583 6598 7584
rect 7754 7648 8070 7649
rect 7754 7584 7760 7648
rect 7824 7584 7840 7648
rect 7904 7584 7920 7648
rect 7984 7584 8000 7648
rect 8064 7584 8070 7648
rect 7754 7583 8070 7584
rect 2602 7104 2918 7105
rect 2602 7040 2608 7104
rect 2672 7040 2688 7104
rect 2752 7040 2768 7104
rect 2832 7040 2848 7104
rect 2912 7040 2918 7104
rect 2602 7039 2918 7040
rect 4074 7104 4390 7105
rect 4074 7040 4080 7104
rect 4144 7040 4160 7104
rect 4224 7040 4240 7104
rect 4304 7040 4320 7104
rect 4384 7040 4390 7104
rect 4074 7039 4390 7040
rect 5546 7104 5862 7105
rect 5546 7040 5552 7104
rect 5616 7040 5632 7104
rect 5696 7040 5712 7104
rect 5776 7040 5792 7104
rect 5856 7040 5862 7104
rect 5546 7039 5862 7040
rect 7018 7104 7334 7105
rect 7018 7040 7024 7104
rect 7088 7040 7104 7104
rect 7168 7040 7184 7104
rect 7248 7040 7264 7104
rect 7328 7040 7334 7104
rect 7018 7039 7334 7040
rect 3338 6560 3654 6561
rect 3338 6496 3344 6560
rect 3408 6496 3424 6560
rect 3488 6496 3504 6560
rect 3568 6496 3584 6560
rect 3648 6496 3654 6560
rect 3338 6495 3654 6496
rect 4810 6560 5126 6561
rect 4810 6496 4816 6560
rect 4880 6496 4896 6560
rect 4960 6496 4976 6560
rect 5040 6496 5056 6560
rect 5120 6496 5126 6560
rect 4810 6495 5126 6496
rect 6282 6560 6598 6561
rect 6282 6496 6288 6560
rect 6352 6496 6368 6560
rect 6432 6496 6448 6560
rect 6512 6496 6528 6560
rect 6592 6496 6598 6560
rect 6282 6495 6598 6496
rect 7754 6560 8070 6561
rect 7754 6496 7760 6560
rect 7824 6496 7840 6560
rect 7904 6496 7920 6560
rect 7984 6496 8000 6560
rect 8064 6496 8070 6560
rect 7754 6495 8070 6496
rect 7465 6082 7531 6085
rect 9600 6082 10000 6112
rect 7465 6080 10000 6082
rect 7465 6024 7470 6080
rect 7526 6024 10000 6080
rect 7465 6022 10000 6024
rect 7465 6019 7531 6022
rect 2602 6016 2918 6017
rect 2602 5952 2608 6016
rect 2672 5952 2688 6016
rect 2752 5952 2768 6016
rect 2832 5952 2848 6016
rect 2912 5952 2918 6016
rect 2602 5951 2918 5952
rect 4074 6016 4390 6017
rect 4074 5952 4080 6016
rect 4144 5952 4160 6016
rect 4224 5952 4240 6016
rect 4304 5952 4320 6016
rect 4384 5952 4390 6016
rect 4074 5951 4390 5952
rect 5546 6016 5862 6017
rect 5546 5952 5552 6016
rect 5616 5952 5632 6016
rect 5696 5952 5712 6016
rect 5776 5952 5792 6016
rect 5856 5952 5862 6016
rect 5546 5951 5862 5952
rect 7018 6016 7334 6017
rect 7018 5952 7024 6016
rect 7088 5952 7104 6016
rect 7168 5952 7184 6016
rect 7248 5952 7264 6016
rect 7328 5952 7334 6016
rect 9600 5992 10000 6022
rect 7018 5951 7334 5952
rect 3338 5472 3654 5473
rect 3338 5408 3344 5472
rect 3408 5408 3424 5472
rect 3488 5408 3504 5472
rect 3568 5408 3584 5472
rect 3648 5408 3654 5472
rect 3338 5407 3654 5408
rect 4810 5472 5126 5473
rect 4810 5408 4816 5472
rect 4880 5408 4896 5472
rect 4960 5408 4976 5472
rect 5040 5408 5056 5472
rect 5120 5408 5126 5472
rect 4810 5407 5126 5408
rect 6282 5472 6598 5473
rect 6282 5408 6288 5472
rect 6352 5408 6368 5472
rect 6432 5408 6448 5472
rect 6512 5408 6528 5472
rect 6592 5408 6598 5472
rect 6282 5407 6598 5408
rect 7754 5472 8070 5473
rect 7754 5408 7760 5472
rect 7824 5408 7840 5472
rect 7904 5408 7920 5472
rect 7984 5408 8000 5472
rect 8064 5408 8070 5472
rect 7754 5407 8070 5408
rect 2602 4928 2918 4929
rect 2602 4864 2608 4928
rect 2672 4864 2688 4928
rect 2752 4864 2768 4928
rect 2832 4864 2848 4928
rect 2912 4864 2918 4928
rect 2602 4863 2918 4864
rect 4074 4928 4390 4929
rect 4074 4864 4080 4928
rect 4144 4864 4160 4928
rect 4224 4864 4240 4928
rect 4304 4864 4320 4928
rect 4384 4864 4390 4928
rect 4074 4863 4390 4864
rect 5546 4928 5862 4929
rect 5546 4864 5552 4928
rect 5616 4864 5632 4928
rect 5696 4864 5712 4928
rect 5776 4864 5792 4928
rect 5856 4864 5862 4928
rect 5546 4863 5862 4864
rect 7018 4928 7334 4929
rect 7018 4864 7024 4928
rect 7088 4864 7104 4928
rect 7168 4864 7184 4928
rect 7248 4864 7264 4928
rect 7328 4864 7334 4928
rect 7018 4863 7334 4864
rect 3338 4384 3654 4385
rect 3338 4320 3344 4384
rect 3408 4320 3424 4384
rect 3488 4320 3504 4384
rect 3568 4320 3584 4384
rect 3648 4320 3654 4384
rect 3338 4319 3654 4320
rect 4810 4384 5126 4385
rect 4810 4320 4816 4384
rect 4880 4320 4896 4384
rect 4960 4320 4976 4384
rect 5040 4320 5056 4384
rect 5120 4320 5126 4384
rect 4810 4319 5126 4320
rect 6282 4384 6598 4385
rect 6282 4320 6288 4384
rect 6352 4320 6368 4384
rect 6432 4320 6448 4384
rect 6512 4320 6528 4384
rect 6592 4320 6598 4384
rect 6282 4319 6598 4320
rect 7754 4384 8070 4385
rect 7754 4320 7760 4384
rect 7824 4320 7840 4384
rect 7904 4320 7920 4384
rect 7984 4320 8000 4384
rect 8064 4320 8070 4384
rect 7754 4319 8070 4320
rect 2602 3840 2918 3841
rect 2602 3776 2608 3840
rect 2672 3776 2688 3840
rect 2752 3776 2768 3840
rect 2832 3776 2848 3840
rect 2912 3776 2918 3840
rect 2602 3775 2918 3776
rect 4074 3840 4390 3841
rect 4074 3776 4080 3840
rect 4144 3776 4160 3840
rect 4224 3776 4240 3840
rect 4304 3776 4320 3840
rect 4384 3776 4390 3840
rect 4074 3775 4390 3776
rect 5546 3840 5862 3841
rect 5546 3776 5552 3840
rect 5616 3776 5632 3840
rect 5696 3776 5712 3840
rect 5776 3776 5792 3840
rect 5856 3776 5862 3840
rect 5546 3775 5862 3776
rect 7018 3840 7334 3841
rect 7018 3776 7024 3840
rect 7088 3776 7104 3840
rect 7168 3776 7184 3840
rect 7248 3776 7264 3840
rect 7328 3776 7334 3840
rect 7018 3775 7334 3776
rect 3338 3296 3654 3297
rect 3338 3232 3344 3296
rect 3408 3232 3424 3296
rect 3488 3232 3504 3296
rect 3568 3232 3584 3296
rect 3648 3232 3654 3296
rect 3338 3231 3654 3232
rect 4810 3296 5126 3297
rect 4810 3232 4816 3296
rect 4880 3232 4896 3296
rect 4960 3232 4976 3296
rect 5040 3232 5056 3296
rect 5120 3232 5126 3296
rect 4810 3231 5126 3232
rect 6282 3296 6598 3297
rect 6282 3232 6288 3296
rect 6352 3232 6368 3296
rect 6432 3232 6448 3296
rect 6512 3232 6528 3296
rect 6592 3232 6598 3296
rect 6282 3231 6598 3232
rect 7754 3296 8070 3297
rect 7754 3232 7760 3296
rect 7824 3232 7840 3296
rect 7904 3232 7920 3296
rect 7984 3232 8000 3296
rect 8064 3232 8070 3296
rect 7754 3231 8070 3232
rect 2602 2752 2918 2753
rect 2602 2688 2608 2752
rect 2672 2688 2688 2752
rect 2752 2688 2768 2752
rect 2832 2688 2848 2752
rect 2912 2688 2918 2752
rect 2602 2687 2918 2688
rect 4074 2752 4390 2753
rect 4074 2688 4080 2752
rect 4144 2688 4160 2752
rect 4224 2688 4240 2752
rect 4304 2688 4320 2752
rect 4384 2688 4390 2752
rect 4074 2687 4390 2688
rect 5546 2752 5862 2753
rect 5546 2688 5552 2752
rect 5616 2688 5632 2752
rect 5696 2688 5712 2752
rect 5776 2688 5792 2752
rect 5856 2688 5862 2752
rect 5546 2687 5862 2688
rect 7018 2752 7334 2753
rect 7018 2688 7024 2752
rect 7088 2688 7104 2752
rect 7168 2688 7184 2752
rect 7248 2688 7264 2752
rect 7328 2688 7334 2752
rect 7018 2687 7334 2688
rect 8201 2274 8267 2277
rect 9600 2274 10000 2304
rect 8201 2272 10000 2274
rect 8201 2216 8206 2272
rect 8262 2216 10000 2272
rect 8201 2214 10000 2216
rect 8201 2211 8267 2214
rect 3338 2208 3654 2209
rect 3338 2144 3344 2208
rect 3408 2144 3424 2208
rect 3488 2144 3504 2208
rect 3568 2144 3584 2208
rect 3648 2144 3654 2208
rect 3338 2143 3654 2144
rect 4810 2208 5126 2209
rect 4810 2144 4816 2208
rect 4880 2144 4896 2208
rect 4960 2144 4976 2208
rect 5040 2144 5056 2208
rect 5120 2144 5126 2208
rect 4810 2143 5126 2144
rect 6282 2208 6598 2209
rect 6282 2144 6288 2208
rect 6352 2144 6368 2208
rect 6432 2144 6448 2208
rect 6512 2144 6528 2208
rect 6592 2144 6598 2208
rect 6282 2143 6598 2144
rect 7754 2208 8070 2209
rect 7754 2144 7760 2208
rect 7824 2144 7840 2208
rect 7904 2144 7920 2208
rect 7984 2144 8000 2208
rect 8064 2144 8070 2208
rect 9600 2184 10000 2214
rect 7754 2143 8070 2144
<< via3 >>
rect 2608 13628 2672 13632
rect 2608 13572 2612 13628
rect 2612 13572 2668 13628
rect 2668 13572 2672 13628
rect 2608 13568 2672 13572
rect 2688 13628 2752 13632
rect 2688 13572 2692 13628
rect 2692 13572 2748 13628
rect 2748 13572 2752 13628
rect 2688 13568 2752 13572
rect 2768 13628 2832 13632
rect 2768 13572 2772 13628
rect 2772 13572 2828 13628
rect 2828 13572 2832 13628
rect 2768 13568 2832 13572
rect 2848 13628 2912 13632
rect 2848 13572 2852 13628
rect 2852 13572 2908 13628
rect 2908 13572 2912 13628
rect 2848 13568 2912 13572
rect 4080 13628 4144 13632
rect 4080 13572 4084 13628
rect 4084 13572 4140 13628
rect 4140 13572 4144 13628
rect 4080 13568 4144 13572
rect 4160 13628 4224 13632
rect 4160 13572 4164 13628
rect 4164 13572 4220 13628
rect 4220 13572 4224 13628
rect 4160 13568 4224 13572
rect 4240 13628 4304 13632
rect 4240 13572 4244 13628
rect 4244 13572 4300 13628
rect 4300 13572 4304 13628
rect 4240 13568 4304 13572
rect 4320 13628 4384 13632
rect 4320 13572 4324 13628
rect 4324 13572 4380 13628
rect 4380 13572 4384 13628
rect 4320 13568 4384 13572
rect 5552 13628 5616 13632
rect 5552 13572 5556 13628
rect 5556 13572 5612 13628
rect 5612 13572 5616 13628
rect 5552 13568 5616 13572
rect 5632 13628 5696 13632
rect 5632 13572 5636 13628
rect 5636 13572 5692 13628
rect 5692 13572 5696 13628
rect 5632 13568 5696 13572
rect 5712 13628 5776 13632
rect 5712 13572 5716 13628
rect 5716 13572 5772 13628
rect 5772 13572 5776 13628
rect 5712 13568 5776 13572
rect 5792 13628 5856 13632
rect 5792 13572 5796 13628
rect 5796 13572 5852 13628
rect 5852 13572 5856 13628
rect 5792 13568 5856 13572
rect 7024 13628 7088 13632
rect 7024 13572 7028 13628
rect 7028 13572 7084 13628
rect 7084 13572 7088 13628
rect 7024 13568 7088 13572
rect 7104 13628 7168 13632
rect 7104 13572 7108 13628
rect 7108 13572 7164 13628
rect 7164 13572 7168 13628
rect 7104 13568 7168 13572
rect 7184 13628 7248 13632
rect 7184 13572 7188 13628
rect 7188 13572 7244 13628
rect 7244 13572 7248 13628
rect 7184 13568 7248 13572
rect 7264 13628 7328 13632
rect 7264 13572 7268 13628
rect 7268 13572 7324 13628
rect 7324 13572 7328 13628
rect 7264 13568 7328 13572
rect 3344 13084 3408 13088
rect 3344 13028 3348 13084
rect 3348 13028 3404 13084
rect 3404 13028 3408 13084
rect 3344 13024 3408 13028
rect 3424 13084 3488 13088
rect 3424 13028 3428 13084
rect 3428 13028 3484 13084
rect 3484 13028 3488 13084
rect 3424 13024 3488 13028
rect 3504 13084 3568 13088
rect 3504 13028 3508 13084
rect 3508 13028 3564 13084
rect 3564 13028 3568 13084
rect 3504 13024 3568 13028
rect 3584 13084 3648 13088
rect 3584 13028 3588 13084
rect 3588 13028 3644 13084
rect 3644 13028 3648 13084
rect 3584 13024 3648 13028
rect 4816 13084 4880 13088
rect 4816 13028 4820 13084
rect 4820 13028 4876 13084
rect 4876 13028 4880 13084
rect 4816 13024 4880 13028
rect 4896 13084 4960 13088
rect 4896 13028 4900 13084
rect 4900 13028 4956 13084
rect 4956 13028 4960 13084
rect 4896 13024 4960 13028
rect 4976 13084 5040 13088
rect 4976 13028 4980 13084
rect 4980 13028 5036 13084
rect 5036 13028 5040 13084
rect 4976 13024 5040 13028
rect 5056 13084 5120 13088
rect 5056 13028 5060 13084
rect 5060 13028 5116 13084
rect 5116 13028 5120 13084
rect 5056 13024 5120 13028
rect 6288 13084 6352 13088
rect 6288 13028 6292 13084
rect 6292 13028 6348 13084
rect 6348 13028 6352 13084
rect 6288 13024 6352 13028
rect 6368 13084 6432 13088
rect 6368 13028 6372 13084
rect 6372 13028 6428 13084
rect 6428 13028 6432 13084
rect 6368 13024 6432 13028
rect 6448 13084 6512 13088
rect 6448 13028 6452 13084
rect 6452 13028 6508 13084
rect 6508 13028 6512 13084
rect 6448 13024 6512 13028
rect 6528 13084 6592 13088
rect 6528 13028 6532 13084
rect 6532 13028 6588 13084
rect 6588 13028 6592 13084
rect 6528 13024 6592 13028
rect 7760 13084 7824 13088
rect 7760 13028 7764 13084
rect 7764 13028 7820 13084
rect 7820 13028 7824 13084
rect 7760 13024 7824 13028
rect 7840 13084 7904 13088
rect 7840 13028 7844 13084
rect 7844 13028 7900 13084
rect 7900 13028 7904 13084
rect 7840 13024 7904 13028
rect 7920 13084 7984 13088
rect 7920 13028 7924 13084
rect 7924 13028 7980 13084
rect 7980 13028 7984 13084
rect 7920 13024 7984 13028
rect 8000 13084 8064 13088
rect 8000 13028 8004 13084
rect 8004 13028 8060 13084
rect 8060 13028 8064 13084
rect 8000 13024 8064 13028
rect 2608 12540 2672 12544
rect 2608 12484 2612 12540
rect 2612 12484 2668 12540
rect 2668 12484 2672 12540
rect 2608 12480 2672 12484
rect 2688 12540 2752 12544
rect 2688 12484 2692 12540
rect 2692 12484 2748 12540
rect 2748 12484 2752 12540
rect 2688 12480 2752 12484
rect 2768 12540 2832 12544
rect 2768 12484 2772 12540
rect 2772 12484 2828 12540
rect 2828 12484 2832 12540
rect 2768 12480 2832 12484
rect 2848 12540 2912 12544
rect 2848 12484 2852 12540
rect 2852 12484 2908 12540
rect 2908 12484 2912 12540
rect 2848 12480 2912 12484
rect 4080 12540 4144 12544
rect 4080 12484 4084 12540
rect 4084 12484 4140 12540
rect 4140 12484 4144 12540
rect 4080 12480 4144 12484
rect 4160 12540 4224 12544
rect 4160 12484 4164 12540
rect 4164 12484 4220 12540
rect 4220 12484 4224 12540
rect 4160 12480 4224 12484
rect 4240 12540 4304 12544
rect 4240 12484 4244 12540
rect 4244 12484 4300 12540
rect 4300 12484 4304 12540
rect 4240 12480 4304 12484
rect 4320 12540 4384 12544
rect 4320 12484 4324 12540
rect 4324 12484 4380 12540
rect 4380 12484 4384 12540
rect 4320 12480 4384 12484
rect 5552 12540 5616 12544
rect 5552 12484 5556 12540
rect 5556 12484 5612 12540
rect 5612 12484 5616 12540
rect 5552 12480 5616 12484
rect 5632 12540 5696 12544
rect 5632 12484 5636 12540
rect 5636 12484 5692 12540
rect 5692 12484 5696 12540
rect 5632 12480 5696 12484
rect 5712 12540 5776 12544
rect 5712 12484 5716 12540
rect 5716 12484 5772 12540
rect 5772 12484 5776 12540
rect 5712 12480 5776 12484
rect 5792 12540 5856 12544
rect 5792 12484 5796 12540
rect 5796 12484 5852 12540
rect 5852 12484 5856 12540
rect 5792 12480 5856 12484
rect 7024 12540 7088 12544
rect 7024 12484 7028 12540
rect 7028 12484 7084 12540
rect 7084 12484 7088 12540
rect 7024 12480 7088 12484
rect 7104 12540 7168 12544
rect 7104 12484 7108 12540
rect 7108 12484 7164 12540
rect 7164 12484 7168 12540
rect 7104 12480 7168 12484
rect 7184 12540 7248 12544
rect 7184 12484 7188 12540
rect 7188 12484 7244 12540
rect 7244 12484 7248 12540
rect 7184 12480 7248 12484
rect 7264 12540 7328 12544
rect 7264 12484 7268 12540
rect 7268 12484 7324 12540
rect 7324 12484 7328 12540
rect 7264 12480 7328 12484
rect 3344 11996 3408 12000
rect 3344 11940 3348 11996
rect 3348 11940 3404 11996
rect 3404 11940 3408 11996
rect 3344 11936 3408 11940
rect 3424 11996 3488 12000
rect 3424 11940 3428 11996
rect 3428 11940 3484 11996
rect 3484 11940 3488 11996
rect 3424 11936 3488 11940
rect 3504 11996 3568 12000
rect 3504 11940 3508 11996
rect 3508 11940 3564 11996
rect 3564 11940 3568 11996
rect 3504 11936 3568 11940
rect 3584 11996 3648 12000
rect 3584 11940 3588 11996
rect 3588 11940 3644 11996
rect 3644 11940 3648 11996
rect 3584 11936 3648 11940
rect 4816 11996 4880 12000
rect 4816 11940 4820 11996
rect 4820 11940 4876 11996
rect 4876 11940 4880 11996
rect 4816 11936 4880 11940
rect 4896 11996 4960 12000
rect 4896 11940 4900 11996
rect 4900 11940 4956 11996
rect 4956 11940 4960 11996
rect 4896 11936 4960 11940
rect 4976 11996 5040 12000
rect 4976 11940 4980 11996
rect 4980 11940 5036 11996
rect 5036 11940 5040 11996
rect 4976 11936 5040 11940
rect 5056 11996 5120 12000
rect 5056 11940 5060 11996
rect 5060 11940 5116 11996
rect 5116 11940 5120 11996
rect 5056 11936 5120 11940
rect 6288 11996 6352 12000
rect 6288 11940 6292 11996
rect 6292 11940 6348 11996
rect 6348 11940 6352 11996
rect 6288 11936 6352 11940
rect 6368 11996 6432 12000
rect 6368 11940 6372 11996
rect 6372 11940 6428 11996
rect 6428 11940 6432 11996
rect 6368 11936 6432 11940
rect 6448 11996 6512 12000
rect 6448 11940 6452 11996
rect 6452 11940 6508 11996
rect 6508 11940 6512 11996
rect 6448 11936 6512 11940
rect 6528 11996 6592 12000
rect 6528 11940 6532 11996
rect 6532 11940 6588 11996
rect 6588 11940 6592 11996
rect 6528 11936 6592 11940
rect 7760 11996 7824 12000
rect 7760 11940 7764 11996
rect 7764 11940 7820 11996
rect 7820 11940 7824 11996
rect 7760 11936 7824 11940
rect 7840 11996 7904 12000
rect 7840 11940 7844 11996
rect 7844 11940 7900 11996
rect 7900 11940 7904 11996
rect 7840 11936 7904 11940
rect 7920 11996 7984 12000
rect 7920 11940 7924 11996
rect 7924 11940 7980 11996
rect 7980 11940 7984 11996
rect 7920 11936 7984 11940
rect 8000 11996 8064 12000
rect 8000 11940 8004 11996
rect 8004 11940 8060 11996
rect 8060 11940 8064 11996
rect 8000 11936 8064 11940
rect 2608 11452 2672 11456
rect 2608 11396 2612 11452
rect 2612 11396 2668 11452
rect 2668 11396 2672 11452
rect 2608 11392 2672 11396
rect 2688 11452 2752 11456
rect 2688 11396 2692 11452
rect 2692 11396 2748 11452
rect 2748 11396 2752 11452
rect 2688 11392 2752 11396
rect 2768 11452 2832 11456
rect 2768 11396 2772 11452
rect 2772 11396 2828 11452
rect 2828 11396 2832 11452
rect 2768 11392 2832 11396
rect 2848 11452 2912 11456
rect 2848 11396 2852 11452
rect 2852 11396 2908 11452
rect 2908 11396 2912 11452
rect 2848 11392 2912 11396
rect 4080 11452 4144 11456
rect 4080 11396 4084 11452
rect 4084 11396 4140 11452
rect 4140 11396 4144 11452
rect 4080 11392 4144 11396
rect 4160 11452 4224 11456
rect 4160 11396 4164 11452
rect 4164 11396 4220 11452
rect 4220 11396 4224 11452
rect 4160 11392 4224 11396
rect 4240 11452 4304 11456
rect 4240 11396 4244 11452
rect 4244 11396 4300 11452
rect 4300 11396 4304 11452
rect 4240 11392 4304 11396
rect 4320 11452 4384 11456
rect 4320 11396 4324 11452
rect 4324 11396 4380 11452
rect 4380 11396 4384 11452
rect 4320 11392 4384 11396
rect 5552 11452 5616 11456
rect 5552 11396 5556 11452
rect 5556 11396 5612 11452
rect 5612 11396 5616 11452
rect 5552 11392 5616 11396
rect 5632 11452 5696 11456
rect 5632 11396 5636 11452
rect 5636 11396 5692 11452
rect 5692 11396 5696 11452
rect 5632 11392 5696 11396
rect 5712 11452 5776 11456
rect 5712 11396 5716 11452
rect 5716 11396 5772 11452
rect 5772 11396 5776 11452
rect 5712 11392 5776 11396
rect 5792 11452 5856 11456
rect 5792 11396 5796 11452
rect 5796 11396 5852 11452
rect 5852 11396 5856 11452
rect 5792 11392 5856 11396
rect 7024 11452 7088 11456
rect 7024 11396 7028 11452
rect 7028 11396 7084 11452
rect 7084 11396 7088 11452
rect 7024 11392 7088 11396
rect 7104 11452 7168 11456
rect 7104 11396 7108 11452
rect 7108 11396 7164 11452
rect 7164 11396 7168 11452
rect 7104 11392 7168 11396
rect 7184 11452 7248 11456
rect 7184 11396 7188 11452
rect 7188 11396 7244 11452
rect 7244 11396 7248 11452
rect 7184 11392 7248 11396
rect 7264 11452 7328 11456
rect 7264 11396 7268 11452
rect 7268 11396 7324 11452
rect 7324 11396 7328 11452
rect 7264 11392 7328 11396
rect 3344 10908 3408 10912
rect 3344 10852 3348 10908
rect 3348 10852 3404 10908
rect 3404 10852 3408 10908
rect 3344 10848 3408 10852
rect 3424 10908 3488 10912
rect 3424 10852 3428 10908
rect 3428 10852 3484 10908
rect 3484 10852 3488 10908
rect 3424 10848 3488 10852
rect 3504 10908 3568 10912
rect 3504 10852 3508 10908
rect 3508 10852 3564 10908
rect 3564 10852 3568 10908
rect 3504 10848 3568 10852
rect 3584 10908 3648 10912
rect 3584 10852 3588 10908
rect 3588 10852 3644 10908
rect 3644 10852 3648 10908
rect 3584 10848 3648 10852
rect 4816 10908 4880 10912
rect 4816 10852 4820 10908
rect 4820 10852 4876 10908
rect 4876 10852 4880 10908
rect 4816 10848 4880 10852
rect 4896 10908 4960 10912
rect 4896 10852 4900 10908
rect 4900 10852 4956 10908
rect 4956 10852 4960 10908
rect 4896 10848 4960 10852
rect 4976 10908 5040 10912
rect 4976 10852 4980 10908
rect 4980 10852 5036 10908
rect 5036 10852 5040 10908
rect 4976 10848 5040 10852
rect 5056 10908 5120 10912
rect 5056 10852 5060 10908
rect 5060 10852 5116 10908
rect 5116 10852 5120 10908
rect 5056 10848 5120 10852
rect 6288 10908 6352 10912
rect 6288 10852 6292 10908
rect 6292 10852 6348 10908
rect 6348 10852 6352 10908
rect 6288 10848 6352 10852
rect 6368 10908 6432 10912
rect 6368 10852 6372 10908
rect 6372 10852 6428 10908
rect 6428 10852 6432 10908
rect 6368 10848 6432 10852
rect 6448 10908 6512 10912
rect 6448 10852 6452 10908
rect 6452 10852 6508 10908
rect 6508 10852 6512 10908
rect 6448 10848 6512 10852
rect 6528 10908 6592 10912
rect 6528 10852 6532 10908
rect 6532 10852 6588 10908
rect 6588 10852 6592 10908
rect 6528 10848 6592 10852
rect 7760 10908 7824 10912
rect 7760 10852 7764 10908
rect 7764 10852 7820 10908
rect 7820 10852 7824 10908
rect 7760 10848 7824 10852
rect 7840 10908 7904 10912
rect 7840 10852 7844 10908
rect 7844 10852 7900 10908
rect 7900 10852 7904 10908
rect 7840 10848 7904 10852
rect 7920 10908 7984 10912
rect 7920 10852 7924 10908
rect 7924 10852 7980 10908
rect 7980 10852 7984 10908
rect 7920 10848 7984 10852
rect 8000 10908 8064 10912
rect 8000 10852 8004 10908
rect 8004 10852 8060 10908
rect 8060 10852 8064 10908
rect 8000 10848 8064 10852
rect 2608 10364 2672 10368
rect 2608 10308 2612 10364
rect 2612 10308 2668 10364
rect 2668 10308 2672 10364
rect 2608 10304 2672 10308
rect 2688 10364 2752 10368
rect 2688 10308 2692 10364
rect 2692 10308 2748 10364
rect 2748 10308 2752 10364
rect 2688 10304 2752 10308
rect 2768 10364 2832 10368
rect 2768 10308 2772 10364
rect 2772 10308 2828 10364
rect 2828 10308 2832 10364
rect 2768 10304 2832 10308
rect 2848 10364 2912 10368
rect 2848 10308 2852 10364
rect 2852 10308 2908 10364
rect 2908 10308 2912 10364
rect 2848 10304 2912 10308
rect 4080 10364 4144 10368
rect 4080 10308 4084 10364
rect 4084 10308 4140 10364
rect 4140 10308 4144 10364
rect 4080 10304 4144 10308
rect 4160 10364 4224 10368
rect 4160 10308 4164 10364
rect 4164 10308 4220 10364
rect 4220 10308 4224 10364
rect 4160 10304 4224 10308
rect 4240 10364 4304 10368
rect 4240 10308 4244 10364
rect 4244 10308 4300 10364
rect 4300 10308 4304 10364
rect 4240 10304 4304 10308
rect 4320 10364 4384 10368
rect 4320 10308 4324 10364
rect 4324 10308 4380 10364
rect 4380 10308 4384 10364
rect 4320 10304 4384 10308
rect 5552 10364 5616 10368
rect 5552 10308 5556 10364
rect 5556 10308 5612 10364
rect 5612 10308 5616 10364
rect 5552 10304 5616 10308
rect 5632 10364 5696 10368
rect 5632 10308 5636 10364
rect 5636 10308 5692 10364
rect 5692 10308 5696 10364
rect 5632 10304 5696 10308
rect 5712 10364 5776 10368
rect 5712 10308 5716 10364
rect 5716 10308 5772 10364
rect 5772 10308 5776 10364
rect 5712 10304 5776 10308
rect 5792 10364 5856 10368
rect 5792 10308 5796 10364
rect 5796 10308 5852 10364
rect 5852 10308 5856 10364
rect 5792 10304 5856 10308
rect 7024 10364 7088 10368
rect 7024 10308 7028 10364
rect 7028 10308 7084 10364
rect 7084 10308 7088 10364
rect 7024 10304 7088 10308
rect 7104 10364 7168 10368
rect 7104 10308 7108 10364
rect 7108 10308 7164 10364
rect 7164 10308 7168 10364
rect 7104 10304 7168 10308
rect 7184 10364 7248 10368
rect 7184 10308 7188 10364
rect 7188 10308 7244 10364
rect 7244 10308 7248 10364
rect 7184 10304 7248 10308
rect 7264 10364 7328 10368
rect 7264 10308 7268 10364
rect 7268 10308 7324 10364
rect 7324 10308 7328 10364
rect 7264 10304 7328 10308
rect 3344 9820 3408 9824
rect 3344 9764 3348 9820
rect 3348 9764 3404 9820
rect 3404 9764 3408 9820
rect 3344 9760 3408 9764
rect 3424 9820 3488 9824
rect 3424 9764 3428 9820
rect 3428 9764 3484 9820
rect 3484 9764 3488 9820
rect 3424 9760 3488 9764
rect 3504 9820 3568 9824
rect 3504 9764 3508 9820
rect 3508 9764 3564 9820
rect 3564 9764 3568 9820
rect 3504 9760 3568 9764
rect 3584 9820 3648 9824
rect 3584 9764 3588 9820
rect 3588 9764 3644 9820
rect 3644 9764 3648 9820
rect 3584 9760 3648 9764
rect 4816 9820 4880 9824
rect 4816 9764 4820 9820
rect 4820 9764 4876 9820
rect 4876 9764 4880 9820
rect 4816 9760 4880 9764
rect 4896 9820 4960 9824
rect 4896 9764 4900 9820
rect 4900 9764 4956 9820
rect 4956 9764 4960 9820
rect 4896 9760 4960 9764
rect 4976 9820 5040 9824
rect 4976 9764 4980 9820
rect 4980 9764 5036 9820
rect 5036 9764 5040 9820
rect 4976 9760 5040 9764
rect 5056 9820 5120 9824
rect 5056 9764 5060 9820
rect 5060 9764 5116 9820
rect 5116 9764 5120 9820
rect 5056 9760 5120 9764
rect 6288 9820 6352 9824
rect 6288 9764 6292 9820
rect 6292 9764 6348 9820
rect 6348 9764 6352 9820
rect 6288 9760 6352 9764
rect 6368 9820 6432 9824
rect 6368 9764 6372 9820
rect 6372 9764 6428 9820
rect 6428 9764 6432 9820
rect 6368 9760 6432 9764
rect 6448 9820 6512 9824
rect 6448 9764 6452 9820
rect 6452 9764 6508 9820
rect 6508 9764 6512 9820
rect 6448 9760 6512 9764
rect 6528 9820 6592 9824
rect 6528 9764 6532 9820
rect 6532 9764 6588 9820
rect 6588 9764 6592 9820
rect 6528 9760 6592 9764
rect 7760 9820 7824 9824
rect 7760 9764 7764 9820
rect 7764 9764 7820 9820
rect 7820 9764 7824 9820
rect 7760 9760 7824 9764
rect 7840 9820 7904 9824
rect 7840 9764 7844 9820
rect 7844 9764 7900 9820
rect 7900 9764 7904 9820
rect 7840 9760 7904 9764
rect 7920 9820 7984 9824
rect 7920 9764 7924 9820
rect 7924 9764 7980 9820
rect 7980 9764 7984 9820
rect 7920 9760 7984 9764
rect 8000 9820 8064 9824
rect 8000 9764 8004 9820
rect 8004 9764 8060 9820
rect 8060 9764 8064 9820
rect 8000 9760 8064 9764
rect 2608 9276 2672 9280
rect 2608 9220 2612 9276
rect 2612 9220 2668 9276
rect 2668 9220 2672 9276
rect 2608 9216 2672 9220
rect 2688 9276 2752 9280
rect 2688 9220 2692 9276
rect 2692 9220 2748 9276
rect 2748 9220 2752 9276
rect 2688 9216 2752 9220
rect 2768 9276 2832 9280
rect 2768 9220 2772 9276
rect 2772 9220 2828 9276
rect 2828 9220 2832 9276
rect 2768 9216 2832 9220
rect 2848 9276 2912 9280
rect 2848 9220 2852 9276
rect 2852 9220 2908 9276
rect 2908 9220 2912 9276
rect 2848 9216 2912 9220
rect 4080 9276 4144 9280
rect 4080 9220 4084 9276
rect 4084 9220 4140 9276
rect 4140 9220 4144 9276
rect 4080 9216 4144 9220
rect 4160 9276 4224 9280
rect 4160 9220 4164 9276
rect 4164 9220 4220 9276
rect 4220 9220 4224 9276
rect 4160 9216 4224 9220
rect 4240 9276 4304 9280
rect 4240 9220 4244 9276
rect 4244 9220 4300 9276
rect 4300 9220 4304 9276
rect 4240 9216 4304 9220
rect 4320 9276 4384 9280
rect 4320 9220 4324 9276
rect 4324 9220 4380 9276
rect 4380 9220 4384 9276
rect 4320 9216 4384 9220
rect 5552 9276 5616 9280
rect 5552 9220 5556 9276
rect 5556 9220 5612 9276
rect 5612 9220 5616 9276
rect 5552 9216 5616 9220
rect 5632 9276 5696 9280
rect 5632 9220 5636 9276
rect 5636 9220 5692 9276
rect 5692 9220 5696 9276
rect 5632 9216 5696 9220
rect 5712 9276 5776 9280
rect 5712 9220 5716 9276
rect 5716 9220 5772 9276
rect 5772 9220 5776 9276
rect 5712 9216 5776 9220
rect 5792 9276 5856 9280
rect 5792 9220 5796 9276
rect 5796 9220 5852 9276
rect 5852 9220 5856 9276
rect 5792 9216 5856 9220
rect 7024 9276 7088 9280
rect 7024 9220 7028 9276
rect 7028 9220 7084 9276
rect 7084 9220 7088 9276
rect 7024 9216 7088 9220
rect 7104 9276 7168 9280
rect 7104 9220 7108 9276
rect 7108 9220 7164 9276
rect 7164 9220 7168 9276
rect 7104 9216 7168 9220
rect 7184 9276 7248 9280
rect 7184 9220 7188 9276
rect 7188 9220 7244 9276
rect 7244 9220 7248 9276
rect 7184 9216 7248 9220
rect 7264 9276 7328 9280
rect 7264 9220 7268 9276
rect 7268 9220 7324 9276
rect 7324 9220 7328 9276
rect 7264 9216 7328 9220
rect 3344 8732 3408 8736
rect 3344 8676 3348 8732
rect 3348 8676 3404 8732
rect 3404 8676 3408 8732
rect 3344 8672 3408 8676
rect 3424 8732 3488 8736
rect 3424 8676 3428 8732
rect 3428 8676 3484 8732
rect 3484 8676 3488 8732
rect 3424 8672 3488 8676
rect 3504 8732 3568 8736
rect 3504 8676 3508 8732
rect 3508 8676 3564 8732
rect 3564 8676 3568 8732
rect 3504 8672 3568 8676
rect 3584 8732 3648 8736
rect 3584 8676 3588 8732
rect 3588 8676 3644 8732
rect 3644 8676 3648 8732
rect 3584 8672 3648 8676
rect 4816 8732 4880 8736
rect 4816 8676 4820 8732
rect 4820 8676 4876 8732
rect 4876 8676 4880 8732
rect 4816 8672 4880 8676
rect 4896 8732 4960 8736
rect 4896 8676 4900 8732
rect 4900 8676 4956 8732
rect 4956 8676 4960 8732
rect 4896 8672 4960 8676
rect 4976 8732 5040 8736
rect 4976 8676 4980 8732
rect 4980 8676 5036 8732
rect 5036 8676 5040 8732
rect 4976 8672 5040 8676
rect 5056 8732 5120 8736
rect 5056 8676 5060 8732
rect 5060 8676 5116 8732
rect 5116 8676 5120 8732
rect 5056 8672 5120 8676
rect 6288 8732 6352 8736
rect 6288 8676 6292 8732
rect 6292 8676 6348 8732
rect 6348 8676 6352 8732
rect 6288 8672 6352 8676
rect 6368 8732 6432 8736
rect 6368 8676 6372 8732
rect 6372 8676 6428 8732
rect 6428 8676 6432 8732
rect 6368 8672 6432 8676
rect 6448 8732 6512 8736
rect 6448 8676 6452 8732
rect 6452 8676 6508 8732
rect 6508 8676 6512 8732
rect 6448 8672 6512 8676
rect 6528 8732 6592 8736
rect 6528 8676 6532 8732
rect 6532 8676 6588 8732
rect 6588 8676 6592 8732
rect 6528 8672 6592 8676
rect 7760 8732 7824 8736
rect 7760 8676 7764 8732
rect 7764 8676 7820 8732
rect 7820 8676 7824 8732
rect 7760 8672 7824 8676
rect 7840 8732 7904 8736
rect 7840 8676 7844 8732
rect 7844 8676 7900 8732
rect 7900 8676 7904 8732
rect 7840 8672 7904 8676
rect 7920 8732 7984 8736
rect 7920 8676 7924 8732
rect 7924 8676 7980 8732
rect 7980 8676 7984 8732
rect 7920 8672 7984 8676
rect 8000 8732 8064 8736
rect 8000 8676 8004 8732
rect 8004 8676 8060 8732
rect 8060 8676 8064 8732
rect 8000 8672 8064 8676
rect 2608 8188 2672 8192
rect 2608 8132 2612 8188
rect 2612 8132 2668 8188
rect 2668 8132 2672 8188
rect 2608 8128 2672 8132
rect 2688 8188 2752 8192
rect 2688 8132 2692 8188
rect 2692 8132 2748 8188
rect 2748 8132 2752 8188
rect 2688 8128 2752 8132
rect 2768 8188 2832 8192
rect 2768 8132 2772 8188
rect 2772 8132 2828 8188
rect 2828 8132 2832 8188
rect 2768 8128 2832 8132
rect 2848 8188 2912 8192
rect 2848 8132 2852 8188
rect 2852 8132 2908 8188
rect 2908 8132 2912 8188
rect 2848 8128 2912 8132
rect 4080 8188 4144 8192
rect 4080 8132 4084 8188
rect 4084 8132 4140 8188
rect 4140 8132 4144 8188
rect 4080 8128 4144 8132
rect 4160 8188 4224 8192
rect 4160 8132 4164 8188
rect 4164 8132 4220 8188
rect 4220 8132 4224 8188
rect 4160 8128 4224 8132
rect 4240 8188 4304 8192
rect 4240 8132 4244 8188
rect 4244 8132 4300 8188
rect 4300 8132 4304 8188
rect 4240 8128 4304 8132
rect 4320 8188 4384 8192
rect 4320 8132 4324 8188
rect 4324 8132 4380 8188
rect 4380 8132 4384 8188
rect 4320 8128 4384 8132
rect 5552 8188 5616 8192
rect 5552 8132 5556 8188
rect 5556 8132 5612 8188
rect 5612 8132 5616 8188
rect 5552 8128 5616 8132
rect 5632 8188 5696 8192
rect 5632 8132 5636 8188
rect 5636 8132 5692 8188
rect 5692 8132 5696 8188
rect 5632 8128 5696 8132
rect 5712 8188 5776 8192
rect 5712 8132 5716 8188
rect 5716 8132 5772 8188
rect 5772 8132 5776 8188
rect 5712 8128 5776 8132
rect 5792 8188 5856 8192
rect 5792 8132 5796 8188
rect 5796 8132 5852 8188
rect 5852 8132 5856 8188
rect 5792 8128 5856 8132
rect 7024 8188 7088 8192
rect 7024 8132 7028 8188
rect 7028 8132 7084 8188
rect 7084 8132 7088 8188
rect 7024 8128 7088 8132
rect 7104 8188 7168 8192
rect 7104 8132 7108 8188
rect 7108 8132 7164 8188
rect 7164 8132 7168 8188
rect 7104 8128 7168 8132
rect 7184 8188 7248 8192
rect 7184 8132 7188 8188
rect 7188 8132 7244 8188
rect 7244 8132 7248 8188
rect 7184 8128 7248 8132
rect 7264 8188 7328 8192
rect 7264 8132 7268 8188
rect 7268 8132 7324 8188
rect 7324 8132 7328 8188
rect 7264 8128 7328 8132
rect 3344 7644 3408 7648
rect 3344 7588 3348 7644
rect 3348 7588 3404 7644
rect 3404 7588 3408 7644
rect 3344 7584 3408 7588
rect 3424 7644 3488 7648
rect 3424 7588 3428 7644
rect 3428 7588 3484 7644
rect 3484 7588 3488 7644
rect 3424 7584 3488 7588
rect 3504 7644 3568 7648
rect 3504 7588 3508 7644
rect 3508 7588 3564 7644
rect 3564 7588 3568 7644
rect 3504 7584 3568 7588
rect 3584 7644 3648 7648
rect 3584 7588 3588 7644
rect 3588 7588 3644 7644
rect 3644 7588 3648 7644
rect 3584 7584 3648 7588
rect 4816 7644 4880 7648
rect 4816 7588 4820 7644
rect 4820 7588 4876 7644
rect 4876 7588 4880 7644
rect 4816 7584 4880 7588
rect 4896 7644 4960 7648
rect 4896 7588 4900 7644
rect 4900 7588 4956 7644
rect 4956 7588 4960 7644
rect 4896 7584 4960 7588
rect 4976 7644 5040 7648
rect 4976 7588 4980 7644
rect 4980 7588 5036 7644
rect 5036 7588 5040 7644
rect 4976 7584 5040 7588
rect 5056 7644 5120 7648
rect 5056 7588 5060 7644
rect 5060 7588 5116 7644
rect 5116 7588 5120 7644
rect 5056 7584 5120 7588
rect 6288 7644 6352 7648
rect 6288 7588 6292 7644
rect 6292 7588 6348 7644
rect 6348 7588 6352 7644
rect 6288 7584 6352 7588
rect 6368 7644 6432 7648
rect 6368 7588 6372 7644
rect 6372 7588 6428 7644
rect 6428 7588 6432 7644
rect 6368 7584 6432 7588
rect 6448 7644 6512 7648
rect 6448 7588 6452 7644
rect 6452 7588 6508 7644
rect 6508 7588 6512 7644
rect 6448 7584 6512 7588
rect 6528 7644 6592 7648
rect 6528 7588 6532 7644
rect 6532 7588 6588 7644
rect 6588 7588 6592 7644
rect 6528 7584 6592 7588
rect 7760 7644 7824 7648
rect 7760 7588 7764 7644
rect 7764 7588 7820 7644
rect 7820 7588 7824 7644
rect 7760 7584 7824 7588
rect 7840 7644 7904 7648
rect 7840 7588 7844 7644
rect 7844 7588 7900 7644
rect 7900 7588 7904 7644
rect 7840 7584 7904 7588
rect 7920 7644 7984 7648
rect 7920 7588 7924 7644
rect 7924 7588 7980 7644
rect 7980 7588 7984 7644
rect 7920 7584 7984 7588
rect 8000 7644 8064 7648
rect 8000 7588 8004 7644
rect 8004 7588 8060 7644
rect 8060 7588 8064 7644
rect 8000 7584 8064 7588
rect 2608 7100 2672 7104
rect 2608 7044 2612 7100
rect 2612 7044 2668 7100
rect 2668 7044 2672 7100
rect 2608 7040 2672 7044
rect 2688 7100 2752 7104
rect 2688 7044 2692 7100
rect 2692 7044 2748 7100
rect 2748 7044 2752 7100
rect 2688 7040 2752 7044
rect 2768 7100 2832 7104
rect 2768 7044 2772 7100
rect 2772 7044 2828 7100
rect 2828 7044 2832 7100
rect 2768 7040 2832 7044
rect 2848 7100 2912 7104
rect 2848 7044 2852 7100
rect 2852 7044 2908 7100
rect 2908 7044 2912 7100
rect 2848 7040 2912 7044
rect 4080 7100 4144 7104
rect 4080 7044 4084 7100
rect 4084 7044 4140 7100
rect 4140 7044 4144 7100
rect 4080 7040 4144 7044
rect 4160 7100 4224 7104
rect 4160 7044 4164 7100
rect 4164 7044 4220 7100
rect 4220 7044 4224 7100
rect 4160 7040 4224 7044
rect 4240 7100 4304 7104
rect 4240 7044 4244 7100
rect 4244 7044 4300 7100
rect 4300 7044 4304 7100
rect 4240 7040 4304 7044
rect 4320 7100 4384 7104
rect 4320 7044 4324 7100
rect 4324 7044 4380 7100
rect 4380 7044 4384 7100
rect 4320 7040 4384 7044
rect 5552 7100 5616 7104
rect 5552 7044 5556 7100
rect 5556 7044 5612 7100
rect 5612 7044 5616 7100
rect 5552 7040 5616 7044
rect 5632 7100 5696 7104
rect 5632 7044 5636 7100
rect 5636 7044 5692 7100
rect 5692 7044 5696 7100
rect 5632 7040 5696 7044
rect 5712 7100 5776 7104
rect 5712 7044 5716 7100
rect 5716 7044 5772 7100
rect 5772 7044 5776 7100
rect 5712 7040 5776 7044
rect 5792 7100 5856 7104
rect 5792 7044 5796 7100
rect 5796 7044 5852 7100
rect 5852 7044 5856 7100
rect 5792 7040 5856 7044
rect 7024 7100 7088 7104
rect 7024 7044 7028 7100
rect 7028 7044 7084 7100
rect 7084 7044 7088 7100
rect 7024 7040 7088 7044
rect 7104 7100 7168 7104
rect 7104 7044 7108 7100
rect 7108 7044 7164 7100
rect 7164 7044 7168 7100
rect 7104 7040 7168 7044
rect 7184 7100 7248 7104
rect 7184 7044 7188 7100
rect 7188 7044 7244 7100
rect 7244 7044 7248 7100
rect 7184 7040 7248 7044
rect 7264 7100 7328 7104
rect 7264 7044 7268 7100
rect 7268 7044 7324 7100
rect 7324 7044 7328 7100
rect 7264 7040 7328 7044
rect 3344 6556 3408 6560
rect 3344 6500 3348 6556
rect 3348 6500 3404 6556
rect 3404 6500 3408 6556
rect 3344 6496 3408 6500
rect 3424 6556 3488 6560
rect 3424 6500 3428 6556
rect 3428 6500 3484 6556
rect 3484 6500 3488 6556
rect 3424 6496 3488 6500
rect 3504 6556 3568 6560
rect 3504 6500 3508 6556
rect 3508 6500 3564 6556
rect 3564 6500 3568 6556
rect 3504 6496 3568 6500
rect 3584 6556 3648 6560
rect 3584 6500 3588 6556
rect 3588 6500 3644 6556
rect 3644 6500 3648 6556
rect 3584 6496 3648 6500
rect 4816 6556 4880 6560
rect 4816 6500 4820 6556
rect 4820 6500 4876 6556
rect 4876 6500 4880 6556
rect 4816 6496 4880 6500
rect 4896 6556 4960 6560
rect 4896 6500 4900 6556
rect 4900 6500 4956 6556
rect 4956 6500 4960 6556
rect 4896 6496 4960 6500
rect 4976 6556 5040 6560
rect 4976 6500 4980 6556
rect 4980 6500 5036 6556
rect 5036 6500 5040 6556
rect 4976 6496 5040 6500
rect 5056 6556 5120 6560
rect 5056 6500 5060 6556
rect 5060 6500 5116 6556
rect 5116 6500 5120 6556
rect 5056 6496 5120 6500
rect 6288 6556 6352 6560
rect 6288 6500 6292 6556
rect 6292 6500 6348 6556
rect 6348 6500 6352 6556
rect 6288 6496 6352 6500
rect 6368 6556 6432 6560
rect 6368 6500 6372 6556
rect 6372 6500 6428 6556
rect 6428 6500 6432 6556
rect 6368 6496 6432 6500
rect 6448 6556 6512 6560
rect 6448 6500 6452 6556
rect 6452 6500 6508 6556
rect 6508 6500 6512 6556
rect 6448 6496 6512 6500
rect 6528 6556 6592 6560
rect 6528 6500 6532 6556
rect 6532 6500 6588 6556
rect 6588 6500 6592 6556
rect 6528 6496 6592 6500
rect 7760 6556 7824 6560
rect 7760 6500 7764 6556
rect 7764 6500 7820 6556
rect 7820 6500 7824 6556
rect 7760 6496 7824 6500
rect 7840 6556 7904 6560
rect 7840 6500 7844 6556
rect 7844 6500 7900 6556
rect 7900 6500 7904 6556
rect 7840 6496 7904 6500
rect 7920 6556 7984 6560
rect 7920 6500 7924 6556
rect 7924 6500 7980 6556
rect 7980 6500 7984 6556
rect 7920 6496 7984 6500
rect 8000 6556 8064 6560
rect 8000 6500 8004 6556
rect 8004 6500 8060 6556
rect 8060 6500 8064 6556
rect 8000 6496 8064 6500
rect 2608 6012 2672 6016
rect 2608 5956 2612 6012
rect 2612 5956 2668 6012
rect 2668 5956 2672 6012
rect 2608 5952 2672 5956
rect 2688 6012 2752 6016
rect 2688 5956 2692 6012
rect 2692 5956 2748 6012
rect 2748 5956 2752 6012
rect 2688 5952 2752 5956
rect 2768 6012 2832 6016
rect 2768 5956 2772 6012
rect 2772 5956 2828 6012
rect 2828 5956 2832 6012
rect 2768 5952 2832 5956
rect 2848 6012 2912 6016
rect 2848 5956 2852 6012
rect 2852 5956 2908 6012
rect 2908 5956 2912 6012
rect 2848 5952 2912 5956
rect 4080 6012 4144 6016
rect 4080 5956 4084 6012
rect 4084 5956 4140 6012
rect 4140 5956 4144 6012
rect 4080 5952 4144 5956
rect 4160 6012 4224 6016
rect 4160 5956 4164 6012
rect 4164 5956 4220 6012
rect 4220 5956 4224 6012
rect 4160 5952 4224 5956
rect 4240 6012 4304 6016
rect 4240 5956 4244 6012
rect 4244 5956 4300 6012
rect 4300 5956 4304 6012
rect 4240 5952 4304 5956
rect 4320 6012 4384 6016
rect 4320 5956 4324 6012
rect 4324 5956 4380 6012
rect 4380 5956 4384 6012
rect 4320 5952 4384 5956
rect 5552 6012 5616 6016
rect 5552 5956 5556 6012
rect 5556 5956 5612 6012
rect 5612 5956 5616 6012
rect 5552 5952 5616 5956
rect 5632 6012 5696 6016
rect 5632 5956 5636 6012
rect 5636 5956 5692 6012
rect 5692 5956 5696 6012
rect 5632 5952 5696 5956
rect 5712 6012 5776 6016
rect 5712 5956 5716 6012
rect 5716 5956 5772 6012
rect 5772 5956 5776 6012
rect 5712 5952 5776 5956
rect 5792 6012 5856 6016
rect 5792 5956 5796 6012
rect 5796 5956 5852 6012
rect 5852 5956 5856 6012
rect 5792 5952 5856 5956
rect 7024 6012 7088 6016
rect 7024 5956 7028 6012
rect 7028 5956 7084 6012
rect 7084 5956 7088 6012
rect 7024 5952 7088 5956
rect 7104 6012 7168 6016
rect 7104 5956 7108 6012
rect 7108 5956 7164 6012
rect 7164 5956 7168 6012
rect 7104 5952 7168 5956
rect 7184 6012 7248 6016
rect 7184 5956 7188 6012
rect 7188 5956 7244 6012
rect 7244 5956 7248 6012
rect 7184 5952 7248 5956
rect 7264 6012 7328 6016
rect 7264 5956 7268 6012
rect 7268 5956 7324 6012
rect 7324 5956 7328 6012
rect 7264 5952 7328 5956
rect 3344 5468 3408 5472
rect 3344 5412 3348 5468
rect 3348 5412 3404 5468
rect 3404 5412 3408 5468
rect 3344 5408 3408 5412
rect 3424 5468 3488 5472
rect 3424 5412 3428 5468
rect 3428 5412 3484 5468
rect 3484 5412 3488 5468
rect 3424 5408 3488 5412
rect 3504 5468 3568 5472
rect 3504 5412 3508 5468
rect 3508 5412 3564 5468
rect 3564 5412 3568 5468
rect 3504 5408 3568 5412
rect 3584 5468 3648 5472
rect 3584 5412 3588 5468
rect 3588 5412 3644 5468
rect 3644 5412 3648 5468
rect 3584 5408 3648 5412
rect 4816 5468 4880 5472
rect 4816 5412 4820 5468
rect 4820 5412 4876 5468
rect 4876 5412 4880 5468
rect 4816 5408 4880 5412
rect 4896 5468 4960 5472
rect 4896 5412 4900 5468
rect 4900 5412 4956 5468
rect 4956 5412 4960 5468
rect 4896 5408 4960 5412
rect 4976 5468 5040 5472
rect 4976 5412 4980 5468
rect 4980 5412 5036 5468
rect 5036 5412 5040 5468
rect 4976 5408 5040 5412
rect 5056 5468 5120 5472
rect 5056 5412 5060 5468
rect 5060 5412 5116 5468
rect 5116 5412 5120 5468
rect 5056 5408 5120 5412
rect 6288 5468 6352 5472
rect 6288 5412 6292 5468
rect 6292 5412 6348 5468
rect 6348 5412 6352 5468
rect 6288 5408 6352 5412
rect 6368 5468 6432 5472
rect 6368 5412 6372 5468
rect 6372 5412 6428 5468
rect 6428 5412 6432 5468
rect 6368 5408 6432 5412
rect 6448 5468 6512 5472
rect 6448 5412 6452 5468
rect 6452 5412 6508 5468
rect 6508 5412 6512 5468
rect 6448 5408 6512 5412
rect 6528 5468 6592 5472
rect 6528 5412 6532 5468
rect 6532 5412 6588 5468
rect 6588 5412 6592 5468
rect 6528 5408 6592 5412
rect 7760 5468 7824 5472
rect 7760 5412 7764 5468
rect 7764 5412 7820 5468
rect 7820 5412 7824 5468
rect 7760 5408 7824 5412
rect 7840 5468 7904 5472
rect 7840 5412 7844 5468
rect 7844 5412 7900 5468
rect 7900 5412 7904 5468
rect 7840 5408 7904 5412
rect 7920 5468 7984 5472
rect 7920 5412 7924 5468
rect 7924 5412 7980 5468
rect 7980 5412 7984 5468
rect 7920 5408 7984 5412
rect 8000 5468 8064 5472
rect 8000 5412 8004 5468
rect 8004 5412 8060 5468
rect 8060 5412 8064 5468
rect 8000 5408 8064 5412
rect 2608 4924 2672 4928
rect 2608 4868 2612 4924
rect 2612 4868 2668 4924
rect 2668 4868 2672 4924
rect 2608 4864 2672 4868
rect 2688 4924 2752 4928
rect 2688 4868 2692 4924
rect 2692 4868 2748 4924
rect 2748 4868 2752 4924
rect 2688 4864 2752 4868
rect 2768 4924 2832 4928
rect 2768 4868 2772 4924
rect 2772 4868 2828 4924
rect 2828 4868 2832 4924
rect 2768 4864 2832 4868
rect 2848 4924 2912 4928
rect 2848 4868 2852 4924
rect 2852 4868 2908 4924
rect 2908 4868 2912 4924
rect 2848 4864 2912 4868
rect 4080 4924 4144 4928
rect 4080 4868 4084 4924
rect 4084 4868 4140 4924
rect 4140 4868 4144 4924
rect 4080 4864 4144 4868
rect 4160 4924 4224 4928
rect 4160 4868 4164 4924
rect 4164 4868 4220 4924
rect 4220 4868 4224 4924
rect 4160 4864 4224 4868
rect 4240 4924 4304 4928
rect 4240 4868 4244 4924
rect 4244 4868 4300 4924
rect 4300 4868 4304 4924
rect 4240 4864 4304 4868
rect 4320 4924 4384 4928
rect 4320 4868 4324 4924
rect 4324 4868 4380 4924
rect 4380 4868 4384 4924
rect 4320 4864 4384 4868
rect 5552 4924 5616 4928
rect 5552 4868 5556 4924
rect 5556 4868 5612 4924
rect 5612 4868 5616 4924
rect 5552 4864 5616 4868
rect 5632 4924 5696 4928
rect 5632 4868 5636 4924
rect 5636 4868 5692 4924
rect 5692 4868 5696 4924
rect 5632 4864 5696 4868
rect 5712 4924 5776 4928
rect 5712 4868 5716 4924
rect 5716 4868 5772 4924
rect 5772 4868 5776 4924
rect 5712 4864 5776 4868
rect 5792 4924 5856 4928
rect 5792 4868 5796 4924
rect 5796 4868 5852 4924
rect 5852 4868 5856 4924
rect 5792 4864 5856 4868
rect 7024 4924 7088 4928
rect 7024 4868 7028 4924
rect 7028 4868 7084 4924
rect 7084 4868 7088 4924
rect 7024 4864 7088 4868
rect 7104 4924 7168 4928
rect 7104 4868 7108 4924
rect 7108 4868 7164 4924
rect 7164 4868 7168 4924
rect 7104 4864 7168 4868
rect 7184 4924 7248 4928
rect 7184 4868 7188 4924
rect 7188 4868 7244 4924
rect 7244 4868 7248 4924
rect 7184 4864 7248 4868
rect 7264 4924 7328 4928
rect 7264 4868 7268 4924
rect 7268 4868 7324 4924
rect 7324 4868 7328 4924
rect 7264 4864 7328 4868
rect 3344 4380 3408 4384
rect 3344 4324 3348 4380
rect 3348 4324 3404 4380
rect 3404 4324 3408 4380
rect 3344 4320 3408 4324
rect 3424 4380 3488 4384
rect 3424 4324 3428 4380
rect 3428 4324 3484 4380
rect 3484 4324 3488 4380
rect 3424 4320 3488 4324
rect 3504 4380 3568 4384
rect 3504 4324 3508 4380
rect 3508 4324 3564 4380
rect 3564 4324 3568 4380
rect 3504 4320 3568 4324
rect 3584 4380 3648 4384
rect 3584 4324 3588 4380
rect 3588 4324 3644 4380
rect 3644 4324 3648 4380
rect 3584 4320 3648 4324
rect 4816 4380 4880 4384
rect 4816 4324 4820 4380
rect 4820 4324 4876 4380
rect 4876 4324 4880 4380
rect 4816 4320 4880 4324
rect 4896 4380 4960 4384
rect 4896 4324 4900 4380
rect 4900 4324 4956 4380
rect 4956 4324 4960 4380
rect 4896 4320 4960 4324
rect 4976 4380 5040 4384
rect 4976 4324 4980 4380
rect 4980 4324 5036 4380
rect 5036 4324 5040 4380
rect 4976 4320 5040 4324
rect 5056 4380 5120 4384
rect 5056 4324 5060 4380
rect 5060 4324 5116 4380
rect 5116 4324 5120 4380
rect 5056 4320 5120 4324
rect 6288 4380 6352 4384
rect 6288 4324 6292 4380
rect 6292 4324 6348 4380
rect 6348 4324 6352 4380
rect 6288 4320 6352 4324
rect 6368 4380 6432 4384
rect 6368 4324 6372 4380
rect 6372 4324 6428 4380
rect 6428 4324 6432 4380
rect 6368 4320 6432 4324
rect 6448 4380 6512 4384
rect 6448 4324 6452 4380
rect 6452 4324 6508 4380
rect 6508 4324 6512 4380
rect 6448 4320 6512 4324
rect 6528 4380 6592 4384
rect 6528 4324 6532 4380
rect 6532 4324 6588 4380
rect 6588 4324 6592 4380
rect 6528 4320 6592 4324
rect 7760 4380 7824 4384
rect 7760 4324 7764 4380
rect 7764 4324 7820 4380
rect 7820 4324 7824 4380
rect 7760 4320 7824 4324
rect 7840 4380 7904 4384
rect 7840 4324 7844 4380
rect 7844 4324 7900 4380
rect 7900 4324 7904 4380
rect 7840 4320 7904 4324
rect 7920 4380 7984 4384
rect 7920 4324 7924 4380
rect 7924 4324 7980 4380
rect 7980 4324 7984 4380
rect 7920 4320 7984 4324
rect 8000 4380 8064 4384
rect 8000 4324 8004 4380
rect 8004 4324 8060 4380
rect 8060 4324 8064 4380
rect 8000 4320 8064 4324
rect 2608 3836 2672 3840
rect 2608 3780 2612 3836
rect 2612 3780 2668 3836
rect 2668 3780 2672 3836
rect 2608 3776 2672 3780
rect 2688 3836 2752 3840
rect 2688 3780 2692 3836
rect 2692 3780 2748 3836
rect 2748 3780 2752 3836
rect 2688 3776 2752 3780
rect 2768 3836 2832 3840
rect 2768 3780 2772 3836
rect 2772 3780 2828 3836
rect 2828 3780 2832 3836
rect 2768 3776 2832 3780
rect 2848 3836 2912 3840
rect 2848 3780 2852 3836
rect 2852 3780 2908 3836
rect 2908 3780 2912 3836
rect 2848 3776 2912 3780
rect 4080 3836 4144 3840
rect 4080 3780 4084 3836
rect 4084 3780 4140 3836
rect 4140 3780 4144 3836
rect 4080 3776 4144 3780
rect 4160 3836 4224 3840
rect 4160 3780 4164 3836
rect 4164 3780 4220 3836
rect 4220 3780 4224 3836
rect 4160 3776 4224 3780
rect 4240 3836 4304 3840
rect 4240 3780 4244 3836
rect 4244 3780 4300 3836
rect 4300 3780 4304 3836
rect 4240 3776 4304 3780
rect 4320 3836 4384 3840
rect 4320 3780 4324 3836
rect 4324 3780 4380 3836
rect 4380 3780 4384 3836
rect 4320 3776 4384 3780
rect 5552 3836 5616 3840
rect 5552 3780 5556 3836
rect 5556 3780 5612 3836
rect 5612 3780 5616 3836
rect 5552 3776 5616 3780
rect 5632 3836 5696 3840
rect 5632 3780 5636 3836
rect 5636 3780 5692 3836
rect 5692 3780 5696 3836
rect 5632 3776 5696 3780
rect 5712 3836 5776 3840
rect 5712 3780 5716 3836
rect 5716 3780 5772 3836
rect 5772 3780 5776 3836
rect 5712 3776 5776 3780
rect 5792 3836 5856 3840
rect 5792 3780 5796 3836
rect 5796 3780 5852 3836
rect 5852 3780 5856 3836
rect 5792 3776 5856 3780
rect 7024 3836 7088 3840
rect 7024 3780 7028 3836
rect 7028 3780 7084 3836
rect 7084 3780 7088 3836
rect 7024 3776 7088 3780
rect 7104 3836 7168 3840
rect 7104 3780 7108 3836
rect 7108 3780 7164 3836
rect 7164 3780 7168 3836
rect 7104 3776 7168 3780
rect 7184 3836 7248 3840
rect 7184 3780 7188 3836
rect 7188 3780 7244 3836
rect 7244 3780 7248 3836
rect 7184 3776 7248 3780
rect 7264 3836 7328 3840
rect 7264 3780 7268 3836
rect 7268 3780 7324 3836
rect 7324 3780 7328 3836
rect 7264 3776 7328 3780
rect 3344 3292 3408 3296
rect 3344 3236 3348 3292
rect 3348 3236 3404 3292
rect 3404 3236 3408 3292
rect 3344 3232 3408 3236
rect 3424 3292 3488 3296
rect 3424 3236 3428 3292
rect 3428 3236 3484 3292
rect 3484 3236 3488 3292
rect 3424 3232 3488 3236
rect 3504 3292 3568 3296
rect 3504 3236 3508 3292
rect 3508 3236 3564 3292
rect 3564 3236 3568 3292
rect 3504 3232 3568 3236
rect 3584 3292 3648 3296
rect 3584 3236 3588 3292
rect 3588 3236 3644 3292
rect 3644 3236 3648 3292
rect 3584 3232 3648 3236
rect 4816 3292 4880 3296
rect 4816 3236 4820 3292
rect 4820 3236 4876 3292
rect 4876 3236 4880 3292
rect 4816 3232 4880 3236
rect 4896 3292 4960 3296
rect 4896 3236 4900 3292
rect 4900 3236 4956 3292
rect 4956 3236 4960 3292
rect 4896 3232 4960 3236
rect 4976 3292 5040 3296
rect 4976 3236 4980 3292
rect 4980 3236 5036 3292
rect 5036 3236 5040 3292
rect 4976 3232 5040 3236
rect 5056 3292 5120 3296
rect 5056 3236 5060 3292
rect 5060 3236 5116 3292
rect 5116 3236 5120 3292
rect 5056 3232 5120 3236
rect 6288 3292 6352 3296
rect 6288 3236 6292 3292
rect 6292 3236 6348 3292
rect 6348 3236 6352 3292
rect 6288 3232 6352 3236
rect 6368 3292 6432 3296
rect 6368 3236 6372 3292
rect 6372 3236 6428 3292
rect 6428 3236 6432 3292
rect 6368 3232 6432 3236
rect 6448 3292 6512 3296
rect 6448 3236 6452 3292
rect 6452 3236 6508 3292
rect 6508 3236 6512 3292
rect 6448 3232 6512 3236
rect 6528 3292 6592 3296
rect 6528 3236 6532 3292
rect 6532 3236 6588 3292
rect 6588 3236 6592 3292
rect 6528 3232 6592 3236
rect 7760 3292 7824 3296
rect 7760 3236 7764 3292
rect 7764 3236 7820 3292
rect 7820 3236 7824 3292
rect 7760 3232 7824 3236
rect 7840 3292 7904 3296
rect 7840 3236 7844 3292
rect 7844 3236 7900 3292
rect 7900 3236 7904 3292
rect 7840 3232 7904 3236
rect 7920 3292 7984 3296
rect 7920 3236 7924 3292
rect 7924 3236 7980 3292
rect 7980 3236 7984 3292
rect 7920 3232 7984 3236
rect 8000 3292 8064 3296
rect 8000 3236 8004 3292
rect 8004 3236 8060 3292
rect 8060 3236 8064 3292
rect 8000 3232 8064 3236
rect 2608 2748 2672 2752
rect 2608 2692 2612 2748
rect 2612 2692 2668 2748
rect 2668 2692 2672 2748
rect 2608 2688 2672 2692
rect 2688 2748 2752 2752
rect 2688 2692 2692 2748
rect 2692 2692 2748 2748
rect 2748 2692 2752 2748
rect 2688 2688 2752 2692
rect 2768 2748 2832 2752
rect 2768 2692 2772 2748
rect 2772 2692 2828 2748
rect 2828 2692 2832 2748
rect 2768 2688 2832 2692
rect 2848 2748 2912 2752
rect 2848 2692 2852 2748
rect 2852 2692 2908 2748
rect 2908 2692 2912 2748
rect 2848 2688 2912 2692
rect 4080 2748 4144 2752
rect 4080 2692 4084 2748
rect 4084 2692 4140 2748
rect 4140 2692 4144 2748
rect 4080 2688 4144 2692
rect 4160 2748 4224 2752
rect 4160 2692 4164 2748
rect 4164 2692 4220 2748
rect 4220 2692 4224 2748
rect 4160 2688 4224 2692
rect 4240 2748 4304 2752
rect 4240 2692 4244 2748
rect 4244 2692 4300 2748
rect 4300 2692 4304 2748
rect 4240 2688 4304 2692
rect 4320 2748 4384 2752
rect 4320 2692 4324 2748
rect 4324 2692 4380 2748
rect 4380 2692 4384 2748
rect 4320 2688 4384 2692
rect 5552 2748 5616 2752
rect 5552 2692 5556 2748
rect 5556 2692 5612 2748
rect 5612 2692 5616 2748
rect 5552 2688 5616 2692
rect 5632 2748 5696 2752
rect 5632 2692 5636 2748
rect 5636 2692 5692 2748
rect 5692 2692 5696 2748
rect 5632 2688 5696 2692
rect 5712 2748 5776 2752
rect 5712 2692 5716 2748
rect 5716 2692 5772 2748
rect 5772 2692 5776 2748
rect 5712 2688 5776 2692
rect 5792 2748 5856 2752
rect 5792 2692 5796 2748
rect 5796 2692 5852 2748
rect 5852 2692 5856 2748
rect 5792 2688 5856 2692
rect 7024 2748 7088 2752
rect 7024 2692 7028 2748
rect 7028 2692 7084 2748
rect 7084 2692 7088 2748
rect 7024 2688 7088 2692
rect 7104 2748 7168 2752
rect 7104 2692 7108 2748
rect 7108 2692 7164 2748
rect 7164 2692 7168 2748
rect 7104 2688 7168 2692
rect 7184 2748 7248 2752
rect 7184 2692 7188 2748
rect 7188 2692 7244 2748
rect 7244 2692 7248 2748
rect 7184 2688 7248 2692
rect 7264 2748 7328 2752
rect 7264 2692 7268 2748
rect 7268 2692 7324 2748
rect 7324 2692 7328 2748
rect 7264 2688 7328 2692
rect 3344 2204 3408 2208
rect 3344 2148 3348 2204
rect 3348 2148 3404 2204
rect 3404 2148 3408 2204
rect 3344 2144 3408 2148
rect 3424 2204 3488 2208
rect 3424 2148 3428 2204
rect 3428 2148 3484 2204
rect 3484 2148 3488 2204
rect 3424 2144 3488 2148
rect 3504 2204 3568 2208
rect 3504 2148 3508 2204
rect 3508 2148 3564 2204
rect 3564 2148 3568 2204
rect 3504 2144 3568 2148
rect 3584 2204 3648 2208
rect 3584 2148 3588 2204
rect 3588 2148 3644 2204
rect 3644 2148 3648 2204
rect 3584 2144 3648 2148
rect 4816 2204 4880 2208
rect 4816 2148 4820 2204
rect 4820 2148 4876 2204
rect 4876 2148 4880 2204
rect 4816 2144 4880 2148
rect 4896 2204 4960 2208
rect 4896 2148 4900 2204
rect 4900 2148 4956 2204
rect 4956 2148 4960 2204
rect 4896 2144 4960 2148
rect 4976 2204 5040 2208
rect 4976 2148 4980 2204
rect 4980 2148 5036 2204
rect 5036 2148 5040 2204
rect 4976 2144 5040 2148
rect 5056 2204 5120 2208
rect 5056 2148 5060 2204
rect 5060 2148 5116 2204
rect 5116 2148 5120 2204
rect 5056 2144 5120 2148
rect 6288 2204 6352 2208
rect 6288 2148 6292 2204
rect 6292 2148 6348 2204
rect 6348 2148 6352 2204
rect 6288 2144 6352 2148
rect 6368 2204 6432 2208
rect 6368 2148 6372 2204
rect 6372 2148 6428 2204
rect 6428 2148 6432 2204
rect 6368 2144 6432 2148
rect 6448 2204 6512 2208
rect 6448 2148 6452 2204
rect 6452 2148 6508 2204
rect 6508 2148 6512 2204
rect 6448 2144 6512 2148
rect 6528 2204 6592 2208
rect 6528 2148 6532 2204
rect 6532 2148 6588 2204
rect 6588 2148 6592 2204
rect 6528 2144 6592 2148
rect 7760 2204 7824 2208
rect 7760 2148 7764 2204
rect 7764 2148 7820 2204
rect 7820 2148 7824 2204
rect 7760 2144 7824 2148
rect 7840 2204 7904 2208
rect 7840 2148 7844 2204
rect 7844 2148 7900 2204
rect 7900 2148 7904 2204
rect 7840 2144 7904 2148
rect 7920 2204 7984 2208
rect 7920 2148 7924 2204
rect 7924 2148 7980 2204
rect 7980 2148 7984 2204
rect 7920 2144 7984 2148
rect 8000 2204 8064 2208
rect 8000 2148 8004 2204
rect 8004 2148 8060 2204
rect 8060 2148 8064 2204
rect 8000 2144 8064 2148
<< metal4 >>
rect 2600 13632 2920 13648
rect 2600 13568 2608 13632
rect 2672 13568 2688 13632
rect 2752 13568 2768 13632
rect 2832 13568 2848 13632
rect 2912 13568 2920 13632
rect 2600 12544 2920 13568
rect 2600 12480 2608 12544
rect 2672 12480 2688 12544
rect 2752 12480 2768 12544
rect 2832 12480 2848 12544
rect 2912 12480 2920 12544
rect 2600 11456 2920 12480
rect 2600 11392 2608 11456
rect 2672 11392 2688 11456
rect 2752 11392 2768 11456
rect 2832 11392 2848 11456
rect 2912 11392 2920 11456
rect 2600 10368 2920 11392
rect 2600 10304 2608 10368
rect 2672 10304 2688 10368
rect 2752 10304 2768 10368
rect 2832 10304 2848 10368
rect 2912 10304 2920 10368
rect 2600 9280 2920 10304
rect 2600 9216 2608 9280
rect 2672 9216 2688 9280
rect 2752 9216 2768 9280
rect 2832 9216 2848 9280
rect 2912 9216 2920 9280
rect 2600 8192 2920 9216
rect 2600 8128 2608 8192
rect 2672 8128 2688 8192
rect 2752 8128 2768 8192
rect 2832 8128 2848 8192
rect 2912 8128 2920 8192
rect 2600 7104 2920 8128
rect 2600 7040 2608 7104
rect 2672 7040 2688 7104
rect 2752 7040 2768 7104
rect 2832 7040 2848 7104
rect 2912 7040 2920 7104
rect 2600 6016 2920 7040
rect 2600 5952 2608 6016
rect 2672 5952 2688 6016
rect 2752 5952 2768 6016
rect 2832 5952 2848 6016
rect 2912 5952 2920 6016
rect 2600 4928 2920 5952
rect 2600 4864 2608 4928
rect 2672 4864 2688 4928
rect 2752 4864 2768 4928
rect 2832 4864 2848 4928
rect 2912 4864 2920 4928
rect 2600 3840 2920 4864
rect 2600 3776 2608 3840
rect 2672 3776 2688 3840
rect 2752 3776 2768 3840
rect 2832 3776 2848 3840
rect 2912 3776 2920 3840
rect 2600 2752 2920 3776
rect 2600 2688 2608 2752
rect 2672 2688 2688 2752
rect 2752 2688 2768 2752
rect 2832 2688 2848 2752
rect 2912 2688 2920 2752
rect 2600 2128 2920 2688
rect 3336 13088 3656 13648
rect 3336 13024 3344 13088
rect 3408 13024 3424 13088
rect 3488 13024 3504 13088
rect 3568 13024 3584 13088
rect 3648 13024 3656 13088
rect 3336 12000 3656 13024
rect 3336 11936 3344 12000
rect 3408 11936 3424 12000
rect 3488 11936 3504 12000
rect 3568 11936 3584 12000
rect 3648 11936 3656 12000
rect 3336 10912 3656 11936
rect 3336 10848 3344 10912
rect 3408 10848 3424 10912
rect 3488 10848 3504 10912
rect 3568 10848 3584 10912
rect 3648 10848 3656 10912
rect 3336 9824 3656 10848
rect 3336 9760 3344 9824
rect 3408 9760 3424 9824
rect 3488 9760 3504 9824
rect 3568 9760 3584 9824
rect 3648 9760 3656 9824
rect 3336 8736 3656 9760
rect 3336 8672 3344 8736
rect 3408 8672 3424 8736
rect 3488 8672 3504 8736
rect 3568 8672 3584 8736
rect 3648 8672 3656 8736
rect 3336 7648 3656 8672
rect 3336 7584 3344 7648
rect 3408 7584 3424 7648
rect 3488 7584 3504 7648
rect 3568 7584 3584 7648
rect 3648 7584 3656 7648
rect 3336 6560 3656 7584
rect 3336 6496 3344 6560
rect 3408 6496 3424 6560
rect 3488 6496 3504 6560
rect 3568 6496 3584 6560
rect 3648 6496 3656 6560
rect 3336 5472 3656 6496
rect 3336 5408 3344 5472
rect 3408 5408 3424 5472
rect 3488 5408 3504 5472
rect 3568 5408 3584 5472
rect 3648 5408 3656 5472
rect 3336 4384 3656 5408
rect 3336 4320 3344 4384
rect 3408 4320 3424 4384
rect 3488 4320 3504 4384
rect 3568 4320 3584 4384
rect 3648 4320 3656 4384
rect 3336 3296 3656 4320
rect 3336 3232 3344 3296
rect 3408 3232 3424 3296
rect 3488 3232 3504 3296
rect 3568 3232 3584 3296
rect 3648 3232 3656 3296
rect 3336 2208 3656 3232
rect 3336 2144 3344 2208
rect 3408 2144 3424 2208
rect 3488 2144 3504 2208
rect 3568 2144 3584 2208
rect 3648 2144 3656 2208
rect 3336 2128 3656 2144
rect 4072 13632 4392 13648
rect 4072 13568 4080 13632
rect 4144 13568 4160 13632
rect 4224 13568 4240 13632
rect 4304 13568 4320 13632
rect 4384 13568 4392 13632
rect 4072 12544 4392 13568
rect 4072 12480 4080 12544
rect 4144 12480 4160 12544
rect 4224 12480 4240 12544
rect 4304 12480 4320 12544
rect 4384 12480 4392 12544
rect 4072 11456 4392 12480
rect 4072 11392 4080 11456
rect 4144 11392 4160 11456
rect 4224 11392 4240 11456
rect 4304 11392 4320 11456
rect 4384 11392 4392 11456
rect 4072 10368 4392 11392
rect 4072 10304 4080 10368
rect 4144 10304 4160 10368
rect 4224 10304 4240 10368
rect 4304 10304 4320 10368
rect 4384 10304 4392 10368
rect 4072 9280 4392 10304
rect 4072 9216 4080 9280
rect 4144 9216 4160 9280
rect 4224 9216 4240 9280
rect 4304 9216 4320 9280
rect 4384 9216 4392 9280
rect 4072 8192 4392 9216
rect 4072 8128 4080 8192
rect 4144 8128 4160 8192
rect 4224 8128 4240 8192
rect 4304 8128 4320 8192
rect 4384 8128 4392 8192
rect 4072 7104 4392 8128
rect 4072 7040 4080 7104
rect 4144 7040 4160 7104
rect 4224 7040 4240 7104
rect 4304 7040 4320 7104
rect 4384 7040 4392 7104
rect 4072 6016 4392 7040
rect 4072 5952 4080 6016
rect 4144 5952 4160 6016
rect 4224 5952 4240 6016
rect 4304 5952 4320 6016
rect 4384 5952 4392 6016
rect 4072 4928 4392 5952
rect 4072 4864 4080 4928
rect 4144 4864 4160 4928
rect 4224 4864 4240 4928
rect 4304 4864 4320 4928
rect 4384 4864 4392 4928
rect 4072 3840 4392 4864
rect 4072 3776 4080 3840
rect 4144 3776 4160 3840
rect 4224 3776 4240 3840
rect 4304 3776 4320 3840
rect 4384 3776 4392 3840
rect 4072 2752 4392 3776
rect 4072 2688 4080 2752
rect 4144 2688 4160 2752
rect 4224 2688 4240 2752
rect 4304 2688 4320 2752
rect 4384 2688 4392 2752
rect 4072 2128 4392 2688
rect 4808 13088 5128 13648
rect 4808 13024 4816 13088
rect 4880 13024 4896 13088
rect 4960 13024 4976 13088
rect 5040 13024 5056 13088
rect 5120 13024 5128 13088
rect 4808 12000 5128 13024
rect 4808 11936 4816 12000
rect 4880 11936 4896 12000
rect 4960 11936 4976 12000
rect 5040 11936 5056 12000
rect 5120 11936 5128 12000
rect 4808 10912 5128 11936
rect 4808 10848 4816 10912
rect 4880 10848 4896 10912
rect 4960 10848 4976 10912
rect 5040 10848 5056 10912
rect 5120 10848 5128 10912
rect 4808 9824 5128 10848
rect 4808 9760 4816 9824
rect 4880 9760 4896 9824
rect 4960 9760 4976 9824
rect 5040 9760 5056 9824
rect 5120 9760 5128 9824
rect 4808 8736 5128 9760
rect 4808 8672 4816 8736
rect 4880 8672 4896 8736
rect 4960 8672 4976 8736
rect 5040 8672 5056 8736
rect 5120 8672 5128 8736
rect 4808 7648 5128 8672
rect 4808 7584 4816 7648
rect 4880 7584 4896 7648
rect 4960 7584 4976 7648
rect 5040 7584 5056 7648
rect 5120 7584 5128 7648
rect 4808 6560 5128 7584
rect 4808 6496 4816 6560
rect 4880 6496 4896 6560
rect 4960 6496 4976 6560
rect 5040 6496 5056 6560
rect 5120 6496 5128 6560
rect 4808 5472 5128 6496
rect 4808 5408 4816 5472
rect 4880 5408 4896 5472
rect 4960 5408 4976 5472
rect 5040 5408 5056 5472
rect 5120 5408 5128 5472
rect 4808 4384 5128 5408
rect 4808 4320 4816 4384
rect 4880 4320 4896 4384
rect 4960 4320 4976 4384
rect 5040 4320 5056 4384
rect 5120 4320 5128 4384
rect 4808 3296 5128 4320
rect 4808 3232 4816 3296
rect 4880 3232 4896 3296
rect 4960 3232 4976 3296
rect 5040 3232 5056 3296
rect 5120 3232 5128 3296
rect 4808 2208 5128 3232
rect 4808 2144 4816 2208
rect 4880 2144 4896 2208
rect 4960 2144 4976 2208
rect 5040 2144 5056 2208
rect 5120 2144 5128 2208
rect 4808 2128 5128 2144
rect 5544 13632 5864 13648
rect 5544 13568 5552 13632
rect 5616 13568 5632 13632
rect 5696 13568 5712 13632
rect 5776 13568 5792 13632
rect 5856 13568 5864 13632
rect 5544 12544 5864 13568
rect 5544 12480 5552 12544
rect 5616 12480 5632 12544
rect 5696 12480 5712 12544
rect 5776 12480 5792 12544
rect 5856 12480 5864 12544
rect 5544 11456 5864 12480
rect 5544 11392 5552 11456
rect 5616 11392 5632 11456
rect 5696 11392 5712 11456
rect 5776 11392 5792 11456
rect 5856 11392 5864 11456
rect 5544 10368 5864 11392
rect 5544 10304 5552 10368
rect 5616 10304 5632 10368
rect 5696 10304 5712 10368
rect 5776 10304 5792 10368
rect 5856 10304 5864 10368
rect 5544 9280 5864 10304
rect 5544 9216 5552 9280
rect 5616 9216 5632 9280
rect 5696 9216 5712 9280
rect 5776 9216 5792 9280
rect 5856 9216 5864 9280
rect 5544 8192 5864 9216
rect 5544 8128 5552 8192
rect 5616 8128 5632 8192
rect 5696 8128 5712 8192
rect 5776 8128 5792 8192
rect 5856 8128 5864 8192
rect 5544 7104 5864 8128
rect 5544 7040 5552 7104
rect 5616 7040 5632 7104
rect 5696 7040 5712 7104
rect 5776 7040 5792 7104
rect 5856 7040 5864 7104
rect 5544 6016 5864 7040
rect 5544 5952 5552 6016
rect 5616 5952 5632 6016
rect 5696 5952 5712 6016
rect 5776 5952 5792 6016
rect 5856 5952 5864 6016
rect 5544 4928 5864 5952
rect 5544 4864 5552 4928
rect 5616 4864 5632 4928
rect 5696 4864 5712 4928
rect 5776 4864 5792 4928
rect 5856 4864 5864 4928
rect 5544 3840 5864 4864
rect 5544 3776 5552 3840
rect 5616 3776 5632 3840
rect 5696 3776 5712 3840
rect 5776 3776 5792 3840
rect 5856 3776 5864 3840
rect 5544 2752 5864 3776
rect 5544 2688 5552 2752
rect 5616 2688 5632 2752
rect 5696 2688 5712 2752
rect 5776 2688 5792 2752
rect 5856 2688 5864 2752
rect 5544 2128 5864 2688
rect 6280 13088 6600 13648
rect 6280 13024 6288 13088
rect 6352 13024 6368 13088
rect 6432 13024 6448 13088
rect 6512 13024 6528 13088
rect 6592 13024 6600 13088
rect 6280 12000 6600 13024
rect 6280 11936 6288 12000
rect 6352 11936 6368 12000
rect 6432 11936 6448 12000
rect 6512 11936 6528 12000
rect 6592 11936 6600 12000
rect 6280 10912 6600 11936
rect 6280 10848 6288 10912
rect 6352 10848 6368 10912
rect 6432 10848 6448 10912
rect 6512 10848 6528 10912
rect 6592 10848 6600 10912
rect 6280 9824 6600 10848
rect 6280 9760 6288 9824
rect 6352 9760 6368 9824
rect 6432 9760 6448 9824
rect 6512 9760 6528 9824
rect 6592 9760 6600 9824
rect 6280 8736 6600 9760
rect 6280 8672 6288 8736
rect 6352 8672 6368 8736
rect 6432 8672 6448 8736
rect 6512 8672 6528 8736
rect 6592 8672 6600 8736
rect 6280 7648 6600 8672
rect 6280 7584 6288 7648
rect 6352 7584 6368 7648
rect 6432 7584 6448 7648
rect 6512 7584 6528 7648
rect 6592 7584 6600 7648
rect 6280 6560 6600 7584
rect 6280 6496 6288 6560
rect 6352 6496 6368 6560
rect 6432 6496 6448 6560
rect 6512 6496 6528 6560
rect 6592 6496 6600 6560
rect 6280 5472 6600 6496
rect 6280 5408 6288 5472
rect 6352 5408 6368 5472
rect 6432 5408 6448 5472
rect 6512 5408 6528 5472
rect 6592 5408 6600 5472
rect 6280 4384 6600 5408
rect 6280 4320 6288 4384
rect 6352 4320 6368 4384
rect 6432 4320 6448 4384
rect 6512 4320 6528 4384
rect 6592 4320 6600 4384
rect 6280 3296 6600 4320
rect 6280 3232 6288 3296
rect 6352 3232 6368 3296
rect 6432 3232 6448 3296
rect 6512 3232 6528 3296
rect 6592 3232 6600 3296
rect 6280 2208 6600 3232
rect 6280 2144 6288 2208
rect 6352 2144 6368 2208
rect 6432 2144 6448 2208
rect 6512 2144 6528 2208
rect 6592 2144 6600 2208
rect 6280 2128 6600 2144
rect 7016 13632 7336 13648
rect 7016 13568 7024 13632
rect 7088 13568 7104 13632
rect 7168 13568 7184 13632
rect 7248 13568 7264 13632
rect 7328 13568 7336 13632
rect 7016 12544 7336 13568
rect 7016 12480 7024 12544
rect 7088 12480 7104 12544
rect 7168 12480 7184 12544
rect 7248 12480 7264 12544
rect 7328 12480 7336 12544
rect 7016 11456 7336 12480
rect 7016 11392 7024 11456
rect 7088 11392 7104 11456
rect 7168 11392 7184 11456
rect 7248 11392 7264 11456
rect 7328 11392 7336 11456
rect 7016 10368 7336 11392
rect 7016 10304 7024 10368
rect 7088 10304 7104 10368
rect 7168 10304 7184 10368
rect 7248 10304 7264 10368
rect 7328 10304 7336 10368
rect 7016 9280 7336 10304
rect 7016 9216 7024 9280
rect 7088 9216 7104 9280
rect 7168 9216 7184 9280
rect 7248 9216 7264 9280
rect 7328 9216 7336 9280
rect 7016 8192 7336 9216
rect 7016 8128 7024 8192
rect 7088 8128 7104 8192
rect 7168 8128 7184 8192
rect 7248 8128 7264 8192
rect 7328 8128 7336 8192
rect 7016 7104 7336 8128
rect 7016 7040 7024 7104
rect 7088 7040 7104 7104
rect 7168 7040 7184 7104
rect 7248 7040 7264 7104
rect 7328 7040 7336 7104
rect 7016 6016 7336 7040
rect 7016 5952 7024 6016
rect 7088 5952 7104 6016
rect 7168 5952 7184 6016
rect 7248 5952 7264 6016
rect 7328 5952 7336 6016
rect 7016 4928 7336 5952
rect 7016 4864 7024 4928
rect 7088 4864 7104 4928
rect 7168 4864 7184 4928
rect 7248 4864 7264 4928
rect 7328 4864 7336 4928
rect 7016 3840 7336 4864
rect 7016 3776 7024 3840
rect 7088 3776 7104 3840
rect 7168 3776 7184 3840
rect 7248 3776 7264 3840
rect 7328 3776 7336 3840
rect 7016 2752 7336 3776
rect 7016 2688 7024 2752
rect 7088 2688 7104 2752
rect 7168 2688 7184 2752
rect 7248 2688 7264 2752
rect 7328 2688 7336 2752
rect 7016 2128 7336 2688
rect 7752 13088 8072 13648
rect 7752 13024 7760 13088
rect 7824 13024 7840 13088
rect 7904 13024 7920 13088
rect 7984 13024 8000 13088
rect 8064 13024 8072 13088
rect 7752 12000 8072 13024
rect 7752 11936 7760 12000
rect 7824 11936 7840 12000
rect 7904 11936 7920 12000
rect 7984 11936 8000 12000
rect 8064 11936 8072 12000
rect 7752 10912 8072 11936
rect 7752 10848 7760 10912
rect 7824 10848 7840 10912
rect 7904 10848 7920 10912
rect 7984 10848 8000 10912
rect 8064 10848 8072 10912
rect 7752 9824 8072 10848
rect 7752 9760 7760 9824
rect 7824 9760 7840 9824
rect 7904 9760 7920 9824
rect 7984 9760 8000 9824
rect 8064 9760 8072 9824
rect 7752 8736 8072 9760
rect 7752 8672 7760 8736
rect 7824 8672 7840 8736
rect 7904 8672 7920 8736
rect 7984 8672 8000 8736
rect 8064 8672 8072 8736
rect 7752 7648 8072 8672
rect 7752 7584 7760 7648
rect 7824 7584 7840 7648
rect 7904 7584 7920 7648
rect 7984 7584 8000 7648
rect 8064 7584 8072 7648
rect 7752 6560 8072 7584
rect 7752 6496 7760 6560
rect 7824 6496 7840 6560
rect 7904 6496 7920 6560
rect 7984 6496 8000 6560
rect 8064 6496 8072 6560
rect 7752 5472 8072 6496
rect 7752 5408 7760 5472
rect 7824 5408 7840 5472
rect 7904 5408 7920 5472
rect 7984 5408 8000 5472
rect 8064 5408 8072 5472
rect 7752 4384 8072 5408
rect 7752 4320 7760 4384
rect 7824 4320 7840 4384
rect 7904 4320 7920 4384
rect 7984 4320 8000 4384
rect 8064 4320 8072 4384
rect 7752 3296 8072 4320
rect 7752 3232 7760 3296
rect 7824 3232 7840 3296
rect 7904 3232 7920 3296
rect 7984 3232 8000 3296
rect 8064 3232 8072 3296
rect 7752 2208 8072 3232
rect 7752 2144 7760 2208
rect 7824 2144 7840 2208
rect 7904 2144 7920 2208
rect 7984 2144 8000 2208
rect 8064 2144 8072 2208
rect 7752 2128 8072 2144
use sky130_fd_sc_hd__nor2_1  _06_
timestamp 1750755022
transform -1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _07_
timestamp 1750755022
transform 1 0 3128 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _08_
timestamp 1750755022
transform -1 0 3956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _09_
timestamp 1750755022
transform 1 0 5520 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _10_
timestamp 1750755022
transform -1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _11_
timestamp 1750755022
transform 1 0 6716 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _12_
timestamp 1750755022
transform 1 0 7268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _13_
timestamp 1750755022
transform -1 0 7452 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _14_
timestamp 1750755022
transform -1 0 6716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _15_
timestamp 1750755022
transform -1 0 7452 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _16_
timestamp 1750755022
transform -1 0 7176 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _17_
timestamp 1750755022
transform 1 0 6900 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _18_
timestamp 1750755022
transform 1 0 7268 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _19_
timestamp 1750755022
transform -1 0 7544 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_9
timestamp 1750755022
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_17
timestamp 1750755022
transform 1 0 3588 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_25
timestamp 1750755022
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1750755022
transform 1 0 4692 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_41
timestamp 1750755022
transform 1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_3
timestamp 1750755022
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_7
timestamp 1750755022
transform 1 0 2668 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_11
timestamp 1750755022
transform 1 0 3036 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_21
timestamp 1750755022
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_33
timestamp 1750755022
transform 1 0 5060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_37
timestamp 1750755022
transform 1 0 5428 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_47
timestamp 1750755022
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_60
timestamp 1750755022
transform 1 0 7544 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1750755022
transform 1 0 2300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1750755022
transform 1 0 3404 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1750755022
transform 1 0 4508 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1750755022
transform 1 0 4692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1750755022
transform 1 0 5796 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_53
timestamp 1750755022
transform 1 0 6900 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_59
timestamp 1750755022
transform 1 0 7452 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1750755022
transform 1 0 2300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1750755022
transform 1 0 3404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1750755022
transform 1 0 4508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1750755022
transform 1 0 5612 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1750755022
transform 1 0 6716 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1750755022
transform 1 0 7084 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_57
timestamp 1750755022
transform 1 0 7268 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1750755022
transform 1 0 2300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1750755022
transform 1 0 3404 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1750755022
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1750755022
transform 1 0 4692 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1750755022
transform 1 0 5796 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_53
timestamp 1750755022
transform 1 0 6900 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1750755022
transform 1 0 2300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1750755022
transform 1 0 3404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1750755022
transform 1 0 4508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1750755022
transform 1 0 5612 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1750755022
transform 1 0 6716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1750755022
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_57
timestamp 1750755022
transform 1 0 7268 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1750755022
transform 1 0 2300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1750755022
transform 1 0 3404 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1750755022
transform 1 0 4508 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1750755022
transform 1 0 4692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1750755022
transform 1 0 5796 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_59
timestamp 1750755022
transform 1 0 7452 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1750755022
transform 1 0 2300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1750755022
transform 1 0 3404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1750755022
transform 1 0 4508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1750755022
transform 1 0 5612 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_51
timestamp 1750755022
transform 1 0 6716 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1750755022
transform 1 0 2300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1750755022
transform 1 0 3404 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1750755022
transform 1 0 4508 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1750755022
transform 1 0 4692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1750755022
transform 1 0 5796 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_53
timestamp 1750755022
transform 1 0 6900 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1750755022
transform 1 0 2300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1750755022
transform 1 0 3404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1750755022
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1750755022
transform 1 0 5612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1750755022
transform 1 0 6716 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1750755022
transform 1 0 7084 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_57
timestamp 1750755022
transform 1 0 7268 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1750755022
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1750755022
transform 1 0 3404 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1750755022
transform 1 0 4508 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1750755022
transform 1 0 4692 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1750755022
transform 1 0 5796 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_53
timestamp 1750755022
transform 1 0 6900 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1750755022
transform 1 0 2300 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1750755022
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1750755022
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1750755022
transform 1 0 5612 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1750755022
transform 1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1750755022
transform 1 0 7084 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_57
timestamp 1750755022
transform 1 0 7268 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1750755022
transform 1 0 2300 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1750755022
transform 1 0 3404 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1750755022
transform 1 0 4508 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1750755022
transform 1 0 4692 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1750755022
transform 1 0 5796 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_53
timestamp 1750755022
transform 1 0 6900 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1750755022
transform 1 0 2300 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1750755022
transform 1 0 3404 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1750755022
transform 1 0 4508 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1750755022
transform 1 0 5612 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1750755022
transform 1 0 6716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1750755022
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1750755022
transform 1 0 2300 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1750755022
transform 1 0 3404 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1750755022
transform 1 0 4508 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1750755022
transform 1 0 4692 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1750755022
transform 1 0 5796 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_59
timestamp 1750755022
transform 1 0 7452 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1750755022
transform 1 0 2300 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1750755022
transform 1 0 3404 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1750755022
transform 1 0 4508 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1750755022
transform 1 0 5612 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1750755022
transform 1 0 6716 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1750755022
transform 1 0 7084 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_60
timestamp 1750755022
transform 1 0 7544 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1750755022
transform 1 0 2300 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1750755022
transform 1 0 3404 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1750755022
transform 1 0 4508 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1750755022
transform 1 0 4692 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1750755022
transform 1 0 5796 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_53
timestamp 1750755022
transform 1 0 6900 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1750755022
transform 1 0 2300 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1750755022
transform 1 0 3404 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1750755022
transform 1 0 4508 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1750755022
transform 1 0 5612 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1750755022
transform 1 0 6716 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1750755022
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_57
timestamp 1750755022
transform 1 0 7268 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1750755022
transform 1 0 2300 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1750755022
transform 1 0 3404 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1750755022
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1750755022
transform 1 0 4692 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1750755022
transform 1 0 5796 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_53
timestamp 1750755022
transform 1 0 6900 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1750755022
transform 1 0 2300 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1750755022
transform 1 0 3404 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1750755022
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1750755022
transform 1 0 5612 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1750755022
transform 1 0 6716 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1750755022
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_60
timestamp 1750755022
transform 1 0 7544 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_3
timestamp 1750755022
transform 1 0 2300 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_10
timestamp 1750755022
transform 1 0 2944 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_22
timestamp 1750755022
transform 1 0 4048 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1750755022
transform 1 0 4692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_41
timestamp 1750755022
transform 1 0 5796 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_49
timestamp 1750755022
transform 1 0 6532 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1750755022
transform -1 0 7636 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1750755022
transform 1 0 2576 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1750755022
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1750755022
transform 1 0 7268 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1750755022
transform 1 0 7268 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output6
timestamp 1750755022
transform -1 0 7176 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output7
timestamp 1750755022
transform -1 0 2852 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output8
timestamp 1750755022
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output9
timestamp 1750755022
transform 1 0 6072 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output10
timestamp 1750755022
transform -1 0 7176 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_21
timestamp 1750755022
transform 1 0 2024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1750755022
transform -1 0 7912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_22
timestamp 1750755022
transform 1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1750755022
transform -1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_23
timestamp 1750755022
transform 1 0 2024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1750755022
transform -1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_24
timestamp 1750755022
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1750755022
transform -1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_25
timestamp 1750755022
transform 1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1750755022
transform -1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_26
timestamp 1750755022
transform 1 0 2024 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1750755022
transform -1 0 7912 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_27
timestamp 1750755022
transform 1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1750755022
transform -1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_28
timestamp 1750755022
transform 1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1750755022
transform -1 0 7912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_29
timestamp 1750755022
transform 1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1750755022
transform -1 0 7912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_30
timestamp 1750755022
transform 1 0 2024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1750755022
transform -1 0 7912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_31
timestamp 1750755022
transform 1 0 2024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1750755022
transform -1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_32
timestamp 1750755022
transform 1 0 2024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1750755022
transform -1 0 7912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_33
timestamp 1750755022
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1750755022
transform -1 0 7912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_34
timestamp 1750755022
transform 1 0 2024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1750755022
transform -1 0 7912 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_35
timestamp 1750755022
transform 1 0 2024 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1750755022
transform -1 0 7912 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_36
timestamp 1750755022
transform 1 0 2024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1750755022
transform -1 0 7912 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_37
timestamp 1750755022
transform 1 0 2024 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1750755022
transform -1 0 7912 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_38
timestamp 1750755022
transform 1 0 2024 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1750755022
transform -1 0 7912 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_39
timestamp 1750755022
transform 1 0 2024 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1750755022
transform -1 0 7912 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_40
timestamp 1750755022
transform 1 0 2024 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1750755022
transform -1 0 7912 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_41
timestamp 1750755022
transform 1 0 2024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1750755022
transform -1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_42
timestamp 1750755022
transform 1 0 4600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_43
timestamp 1750755022
transform 1 0 7176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp 1750755022
transform 1 0 7176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_45
timestamp 1750755022
transform 1 0 4600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_46
timestamp 1750755022
transform 1 0 7176 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_47
timestamp 1750755022
transform 1 0 4600 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_48
timestamp 1750755022
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_49
timestamp 1750755022
transform 1 0 4600 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_50
timestamp 1750755022
transform 1 0 7176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_51
timestamp 1750755022
transform 1 0 4600 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_52
timestamp 1750755022
transform 1 0 7176 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_53
timestamp 1750755022
transform 1 0 4600 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_54
timestamp 1750755022
transform 1 0 7176 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_55
timestamp 1750755022
transform 1 0 4600 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_56
timestamp 1750755022
transform 1 0 7176 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_57
timestamp 1750755022
transform 1 0 4600 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_58
timestamp 1750755022
transform 1 0 7176 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_59
timestamp 1750755022
transform 1 0 4600 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_60
timestamp 1750755022
transform 1 0 7176 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_61
timestamp 1750755022
transform 1 0 4600 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_62
timestamp 1750755022
transform 1 0 7176 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_63
timestamp 1750755022
transform 1 0 4600 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_64
timestamp 1750755022
transform 1 0 7176 0 1 13056
box -38 -48 130 592
<< labels >>
rlabel metal2 s 5048 13056 5048 13056 4 VGND
rlabel metal1 s 4968 13600 4968 13600 4 VPWR
rlabel metal1 s 3680 3026 3680 3026 4 _00_
rlabel metal1 s 6072 3026 6072 3026 4 _01_
rlabel metal1 s 7314 3026 7314 3026 4 _02_
rlabel metal1 s 6578 3026 6578 3026 4 _03_
rlabel metal2 s 6946 6086 6946 6086 4 _04_
rlabel metal2 s 7406 10438 7406 10438 4 _05_
rlabel metal2 s 7498 14494 7498 14494 4 a
rlabel metal1 s 2622 13294 2622 13294 4 b
rlabel metal3 s 8932 2244 8932 2244 4 d[0]
rlabel metal3 s 8564 6052 8564 6052 4 d[1]
rlabel metal3 s 7843 9996 7843 9996 4 d[2]
rlabel metal1 s 7590 13430 7590 13430 4 d[3]
rlabel metal2 s 1242 1350 1242 1350 4 m[0]
rlabel metal2 s 3726 1316 3726 1316 4 m[1]
rlabel metal2 s 6210 1316 6210 1316 4 m[2]
rlabel metal2 s 8694 1350 8694 1350 4 m[3]
rlabel metal1 s 7360 5882 7360 5882 4 net1
rlabel metal1 s 6992 2414 6992 2414 4 net10
rlabel metal1 s 7498 5678 7498 5678 4 net2
rlabel metal1 s 7360 2414 7360 2414 4 net3
rlabel metal1 s 7222 6290 7222 6290 4 net4
rlabel metal1 s 7452 9554 7452 9554 4 net5
rlabel metal2 s 7314 13090 7314 13090 4 net6
rlabel metal1 s 2852 2414 2852 2414 4 net7
rlabel metal2 s 3910 2618 3910 2618 4 net8
rlabel metal1 s 6256 2414 6256 2414 4 net9
flabel metal4 s 7752 2128 8072 13648 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 6280 2128 6600 13648 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4808 2128 5128 13648 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 3336 2128 3656 13648 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7016 2128 7336 13648 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 5544 2128 5864 13648 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 4072 2128 4392 13648 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2600 2128 2920 13648 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 7470 15600 7526 16000 0 FreeSans 280 90 0 0 a
port 3 nsew
flabel metal2 s 2502 15600 2558 16000 0 FreeSans 280 90 0 0 b
port 4 nsew
flabel metal3 s 9600 2184 10000 2304 0 FreeSans 600 0 0 0 d[0]
port 5 nsew
flabel metal3 s 9600 5992 10000 6112 0 FreeSans 600 0 0 0 d[1]
port 6 nsew
flabel metal3 s 9600 9800 10000 9920 0 FreeSans 600 0 0 0 d[2]
port 7 nsew
flabel metal3 s 9600 13608 10000 13728 0 FreeSans 600 0 0 0 d[3]
port 8 nsew
flabel metal2 s 1214 0 1270 400 0 FreeSans 280 90 0 0 m[0]
port 9 nsew
flabel metal2 s 3698 0 3754 400 0 FreeSans 280 90 0 0 m[1]
port 10 nsew
flabel metal2 s 6182 0 6238 400 0 FreeSans 280 90 0 0 m[2]
port 11 nsew
flabel metal2 s 8666 0 8722 400 0 FreeSans 280 90 0 0 m[3]
port 12 nsew
<< properties >>
string FIXED_BBOX 0 0 10000 16000
string GDS_END 204896
string GDS_FILE ../gds/Decoder.gds
string GDS_START 65708
<< end >>
